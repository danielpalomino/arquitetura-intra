LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;
LIBRARY WORK;
USE WORK.INTRA_LIBRARY.ALL;

ENTITY fp IS
	GENERIC (n: INTEGER:= 8)
	PORT (
		clk,reset: IN STD_LOGIC;
		bs_selectors0, bs_selectors1: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		sample0,sample1: IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		predicted_pixel: OUT STD_LOGIC_VECTOR(n+2 DOWNTO 0)
		);
END fp;

ARCHITECTURE behavior OF fp IS

BEGIN




END behavior;
