LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;

ENTITY neighbor_buffer IS
	GENERIC (n: INTEGER:= 8);
	PORT (
		clk,reset		: IN STD_LOGIC;
		enable			: IN STD_LOGIC;
		mux_above		: IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		mux_left			: IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		input_sample	: IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		neighbor_above0: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		neighbor_above1: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		neighbor_above2: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		neighbor_above3: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		neighbor_above4: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		neighbor_left0	: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		neighbor_left1	: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		neighbor_left2	: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		neighbor_left3	: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		neighbor_left4	: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0)
		);
END neighbor_buffer;

ARCHITECTURE behavior OF neighbor_buffer IS

SIGNAL	neighbor0, neighbor1, neighbor2, neighbor3, neighbor4, neighbor5, neighbor6, neighbor7,
			neighbor8, neighbor9, neighbor10,neighbor11,neighbor12,neighbor13,neighbor14,neighbor15,
			neighbor16,neighbor17,neighbor18,neighbor19,neighbor20,neighbor21,neighbor22,neighbor23,
			neighbor24,neighbor25,neighbor26,neighbor27,neighbor28,neighbor29,neighbor30,neighbor31,
			neighbor32,neighbor33,neighbor34,neighbor35,neighbor36,neighbor37,neighbor38,neighbor39,
			neighbor40,neighbor41,neighbor42,neighbor43,neighbor44,neighbor45,neighbor46,neighbor47,
			neighbor48,neighbor49,neighbor50,neighbor51,neighbor52,neighbor53,neighbor54,neighbor55,
			neighbor56,neighbor57,neighbor58,neighbor59,neighbor60,neighbor61,neighbor62,neighbor63,
			neighborDC,
			neighbor64,neighbor65,neighbor66,neighbor67,neighbor68,neighbor69,neighbor70,neighbor71,
			neighbor72,neighbor73,neighbor74,neighbor75,neighbor76,neighbor77,neighbor78,neighbor79,
			neighbor80,neighbor81,neighbor82,neighbor83,neighbor84,neighbor85,neighbor86,neighbor87,
			neighbor88,neighbor89,neighbor90,neighbor91,neighbor92,neighbor93,neighbor94,neighbor95,
			neighbor96, neighbor97, neighbor98, neighbor99, neighbor100,neighbor101,neighbor102,neighbor103,
			neighbor104,neighbor105,neighbor106,neighbor107,neighbor108,neighbor109,neighbor110,neighbor111,
			neighbor112,neighbor113,neighbor114,neighbor115,neighbor116,neighbor117,neighbor118,neighbor119,
			neighbor120,neighbor121,neighbor122,neighbor123,neighbor124,neighbor125,neighbor126,neighbor127
			: STD_LOGIC_VECTOR (n-1 DOWNTO 0);

BEGIN

	PROCESS (clk,reset)
	BEGIN
		IF reset = '1' THEN
			neighbor0 <= (OTHERS=>'0');
			neighbor1 <= (OTHERS=>'0');
			neighbor2 <= (OTHERS=>'0');
			neighbor3 <= (OTHERS=>'0');
			neighbor4 <= (OTHERS=>'0');
			neighbor5 <= (OTHERS=>'0');
			neighbor6 <= (OTHERS=>'0');
			neighbor7 <= (OTHERS=>'0');
			neighbor8 <= (OTHERS=>'0');
			neighbor9 <= (OTHERS=>'0');
			neighbor10 <= (OTHERS=>'0');
			neighbor11 <= (OTHERS=>'0');
			neighbor12 <= (OTHERS=>'0');
			neighbor13 <= (OTHERS=>'0');
			neighbor14 <= (OTHERS=>'0');
			neighbor15 <= (OTHERS=>'0');
			neighbor16 <= (OTHERS=>'0');
			neighbor17 <= (OTHERS=>'0');
			neighbor18 <= (OTHERS=>'0');
			neighbor19 <= (OTHERS=>'0');
			neighbor20 <= (OTHERS=>'0');
			neighbor21 <= (OTHERS=>'0');
			neighbor22 <= (OTHERS=>'0');
			neighbor23 <= (OTHERS=>'0');
			neighbor24 <= (OTHERS=>'0');
			neighbor25 <= (OTHERS=>'0');
			neighbor26 <= (OTHERS=>'0');
			neighbor27 <= (OTHERS=>'0');
			neighbor28 <= (OTHERS=>'0');
			neighbor29 <= (OTHERS=>'0');
			neighbor30 <= (OTHERS=>'0');
			neighbor31 <= (OTHERS=>'0');
			neighbor32 <= (OTHERS=>'0');
			neighbor33 <= (OTHERS=>'0');
			neighbor34 <= (OTHERS=>'0');
			neighbor35 <= (OTHERS=>'0');
			neighbor36 <= (OTHERS=>'0');
			neighbor37 <= (OTHERS=>'0');
			neighbor38 <= (OTHERS=>'0');
			neighbor39 <= (OTHERS=>'0');
			neighbor40 <= (OTHERS=>'0');
			neighbor41 <= (OTHERS=>'0');
			neighbor42 <= (OTHERS=>'0');
			neighbor43 <= (OTHERS=>'0');
			neighbor44 <= (OTHERS=>'0');
			neighbor45 <= (OTHERS=>'0');
			neighbor46 <= (OTHERS=>'0');
			neighbor47 <= (OTHERS=>'0');
			neighbor48 <= (OTHERS=>'0');
			neighbor49 <= (OTHERS=>'0');
			neighbor50 <= (OTHERS=>'0');
			neighbor51 <= (OTHERS=>'0');
			neighbor52 <= (OTHERS=>'0');
			neighbor53 <= (OTHERS=>'0');
			neighbor54 <= (OTHERS=>'0');
			neighbor55 <= (OTHERS=>'0');
			neighbor56 <= (OTHERS=>'0');
			neighbor57 <= (OTHERS=>'0');
			neighbor58 <= (OTHERS=>'0');
			neighbor59 <= (OTHERS=>'0');
			neighbor60 <= (OTHERS=>'0');
			neighbor61 <= (OTHERS=>'0');
			neighbor62 <= (OTHERS=>'0');
			neighbor63 <= (OTHERS=>'0');
			neighborDC <= (OTHERS=>'0');
			neighbor64 <= (OTHERS=>'0');
			neighbor65 <= (OTHERS=>'0');
			neighbor66 <= (OTHERS=>'0');
			neighbor67 <= (OTHERS=>'0');
			neighbor68 <= (OTHERS=>'0');
			neighbor69 <= (OTHERS=>'0');
			neighbor70 <= (OTHERS=>'0');
			neighbor71 <= (OTHERS=>'0');
			neighbor72 <= (OTHERS=>'0');
			neighbor73 <= (OTHERS=>'0');
			neighbor74 <= (OTHERS=>'0');
			neighbor75 <= (OTHERS=>'0');
			neighbor76 <= (OTHERS=>'0');
			neighbor77 <= (OTHERS=>'0');
			neighbor78 <= (OTHERS=>'0');
			neighbor79 <= (OTHERS=>'0');
			neighbor80 <= (OTHERS=>'0');
			neighbor81 <= (OTHERS=>'0');
			neighbor82 <= (OTHERS=>'0');
			neighbor83 <= (OTHERS=>'0');
			neighbor84 <= (OTHERS=>'0');
			neighbor85 <= (OTHERS=>'0');
			neighbor86 <= (OTHERS=>'0');
			neighbor87 <= (OTHERS=>'0');
			neighbor88 <= (OTHERS=>'0');
			neighbor89 <= (OTHERS=>'0');
			neighbor90 <= (OTHERS=>'0');
			neighbor91 <= (OTHERS=>'0');
			neighbor92 <= (OTHERS=>'0');
			neighbor93 <= (OTHERS=>'0');
			neighbor94 <= (OTHERS=>'0');
			neighbor95 <= (OTHERS=>'0');
			neighbor96 <= (OTHERS=>'0');
			neighbor97 <= (OTHERS=>'0');
			neighbor98 <= (OTHERS=>'0');
			neighbor99 <= (OTHERS=>'0');
			neighbor100 <= (OTHERS=>'0');
			neighbor101 <= (OTHERS=>'0');
			neighbor102 <= (OTHERS=>'0');
			neighbor103 <= (OTHERS=>'0');
			neighbor104 <= (OTHERS=>'0');
			neighbor105 <= (OTHERS=>'0');
			neighbor106 <= (OTHERS=>'0');
			neighbor107 <= (OTHERS=>'0');
			neighbor108 <= (OTHERS=>'0');
			neighbor109 <= (OTHERS=>'0');
			neighbor110 <= (OTHERS=>'0');
			neighbor111 <= (OTHERS=>'0');
			neighbor112 <= (OTHERS=>'0');
			neighbor113 <= (OTHERS=>'0');
			neighbor114 <= (OTHERS=>'0');
			neighbor115 <= (OTHERS=>'0');
			neighbor116 <= (OTHERS=>'0');
			neighbor117 <= (OTHERS=>'0');
			neighbor118 <= (OTHERS=>'0');
			neighbor119 <= (OTHERS=>'0');
			neighbor120 <= (OTHERS=>'0');
			neighbor121 <= (OTHERS=>'0');
			neighbor122 <= (OTHERS=>'0');
			neighbor123 <= (OTHERS=>'0');
			neighbor124 <= (OTHERS=>'0');
			neighbor125 <= (OTHERS=>'0');
			neighbor126 <= (OTHERS=>'0');
			neighbor127 <= (OTHERS=>'0');
		ELSIF clk'EVENT AND clk = '1' THEN
			IF enable = '1' THEN
				neighbor0 <= input_sample;
				neighbor1 <= neighbor0;
				neighbor2 <= neighbor1;
				neighbor3 <= neighbor2;
				neighbor4 <= neighbor3;
				neighbor5 <= neighbor4;
				neighbor6 <= neighbor5;
				neighbor7 <= neighbor6;
				neighbor8 <= neighbor7;
				neighbor9 <= neighbor8;
				neighbor10 <= neighbor9;
				neighbor11 <= neighbor10;
				neighbor12 <= neighbor11;
				neighbor13 <= neighbor12;
				neighbor14 <= neighbor13;
				neighbor15 <= neighbor14;
				neighbor16 <= neighbor15;
				neighbor17 <= neighbor16;
				neighbor18 <= neighbor17;
				neighbor19 <= neighbor18;
				neighbor20 <= neighbor19;
				neighbor21 <= neighbor20;
				neighbor22 <= neighbor21;
				neighbor23 <= neighbor22;
				neighbor24 <= neighbor23;
				neighbor25 <= neighbor24;
				neighbor26 <= neighbor25;
				neighbor27 <= neighbor26;
				neighbor28 <= neighbor27;
				neighbor29 <= neighbor28;
				neighbor30 <= neighbor29;
				neighbor31 <= neighbor30;
				neighbor32 <= neighbor31;
				neighbor33 <= neighbor32;
				neighbor34 <= neighbor33;
				neighbor35 <= neighbor34;
				neighbor36 <= neighbor35;
				neighbor37 <= neighbor36;
				neighbor38 <= neighbor37;
				neighbor39 <= neighbor38;
				neighbor40 <= neighbor39;
				neighbor41 <= neighbor40;
				neighbor42 <= neighbor41;
				neighbor43 <= neighbor42;
				neighbor44 <= neighbor43;
				neighbor45 <= neighbor44;
				neighbor46 <= neighbor45;
				neighbor47 <= neighbor46;
				neighbor48 <= neighbor47;
				neighbor49 <= neighbor48;
				neighbor50 <= neighbor49;
				neighbor51 <= neighbor50;
				neighbor52 <= neighbor51;
				neighbor53 <= neighbor52;
				neighbor54 <= neighbor53;
				neighbor55 <= neighbor54;
				neighbor56 <= neighbor55;
				neighbor57 <= neighbor56;
				neighbor58 <= neighbor57;
				neighbor59 <= neighbor58;
				neighbor60 <= neighbor59;
				neighbor61 <= neighbor60;
				neighbor62 <= neighbor61;
				neighbor63 <= neighbor62;
				
				neighborDC <= neighbor63;
				
				neighbor64 <= neighborDC;
				neighbor65 <= neighbor64;
				neighbor66 <= neighbor65;
				neighbor67 <= neighbor66;
				neighbor68 <= neighbor67;
				neighbor69 <= neighbor68;
				neighbor70 <= neighbor69;
				neighbor71 <= neighbor70;
				neighbor72 <= neighbor71;
				neighbor73 <= neighbor72;
				neighbor74 <= neighbor73;
				neighbor75 <= neighbor74;
				neighbor76 <= neighbor75;
				neighbor77 <= neighbor76;
				neighbor78 <= neighbor77;
				neighbor79 <= neighbor78;
				neighbor80 <= neighbor79;
				neighbor81 <= neighbor80;
				neighbor82 <= neighbor81;
				neighbor83 <= neighbor82;
				neighbor84 <= neighbor83;
				neighbor85 <= neighbor84;
				neighbor86 <= neighbor85;
				neighbor87 <= neighbor86;
				neighbor88 <= neighbor87;
				neighbor89 <= neighbor88;
				neighbor90 <= neighbor89;
				neighbor91 <= neighbor90;
				neighbor92 <= neighbor91;
				neighbor93 <= neighbor92;
				neighbor94 <= neighbor93;
				neighbor95 <= neighbor94;
				neighbor96 <= neighbor95;
				neighbor97 <= neighbor96;
				neighbor98 <= neighbor97;
				neighbor99 <= neighbor98;
				neighbor100 <= neighbor99;
				neighbor101 <= neighbor100;
				neighbor102 <= neighbor101;
				neighbor103 <= neighbor102;
				neighbor104 <= neighbor103;
				neighbor105 <= neighbor104;
				neighbor106 <= neighbor105;
				neighbor107 <= neighbor106;
				neighbor108 <= neighbor107;
				neighbor109 <= neighbor108;
				neighbor110 <= neighbor109;
				neighbor111 <= neighbor110;
				neighbor112 <= neighbor111;
				neighbor113 <= neighbor112;
				neighbor114 <= neighbor113;
				neighbor115 <= neighbor114;
				neighbor116 <= neighbor115;
				neighbor117 <= neighbor116;
				neighbor118 <= neighbor117;
				neighbor119 <= neighbor118;
				neighbor120 <= neighbor119;
				neighbor121 <= neighbor120;
				neighbor122 <= neighbor121;
				neighbor123 <= neighbor122;
				neighbor124 <= neighbor123;
				neighbor125 <= neighbor124;
				neighbor126 <= neighbor125;
				neighbor127 <= neighbor126;
			END IF;
		END IF;
	END PROCESS;
	
	WITH mux_above SELECT
	neighbor_above0	<=	neighbor0	WHEN "0000000",
								neighbor1	WHEN "0000001",
								neighbor2	WHEN "0000010",
								neighbor3	WHEN "0000011",
								neighbor4	WHEN "0000100",
								neighbor5	WHEN "0000101",
								neighbor6	WHEN "0000110",
								neighbor7	WHEN "0000111",
								neighbor8	WHEN "0001000",
								neighbor9	WHEN "0001001",
								neighbor10	WHEN "0001010",
								neighbor11	WHEN "0001011",
								neighbor12	WHEN "0001100",
								neighbor13	WHEN "0001101",
								neighbor14	WHEN "0001110",
								neighbor15	WHEN "0001111",
								neighbor16	WHEN "0010000",
								neighbor17	WHEN "0010001",
								neighbor18	WHEN "0010010",
								neighbor19	WHEN "0010011",
								neighbor20	WHEN "0010100",
								neighbor21	WHEN "0010101",
								neighbor22	WHEN "0010110",
								neighbor23	WHEN "0010111",
								neighbor24	WHEN "0011000",
								neighbor25	WHEN "0011001",
								neighbor26	WHEN "0011010",
								neighbor27	WHEN "0011011",
								neighbor28	WHEN "0011100",
								neighbor29	WHEN "0011101",
								neighbor30	WHEN "0011110",
								neighbor31	WHEN "0011111",
								neighbor32	WHEN "0100000",
								neighbor33	WHEN "0100001",
								neighbor34	WHEN "0100010",
								neighbor35	WHEN "0100011",
								neighbor36	WHEN "0100100",
								neighbor37	WHEN "0100101",
								neighbor38	WHEN "0100110",
								neighbor39	WHEN "0100111",
								neighbor40	WHEN "0101000",
								neighbor41	WHEN "0101001",
								neighbor42	WHEN "0101010",
								neighbor43	WHEN "0101011",
								neighbor44	WHEN "0101100",
								neighbor45	WHEN "0101101",
								neighbor46	WHEN "0101110",
								neighbor47	WHEN "0101111",
								neighbor48	WHEN "0110000",
								neighbor49	WHEN "0110001",
								neighbor50	WHEN "0110010",
								neighbor51	WHEN "0110011",
								neighbor52	WHEN "0110100",
								neighbor53	WHEN "0110101",
								neighbor54	WHEN "0110110",
								neighbor55	WHEN "0110111",
								neighbor56	WHEN "0111000",
								neighbor57	WHEN "0111001",
								neighbor58	WHEN "0111010",
								neighbor59	WHEN "0111011",
								neighbor60	WHEN "0111100",
								neighbor61	WHEN "0111101",
								neighbor62	WHEN "0111110",
								neighbor63	WHEN "0111111",
								
								neighborDC	WHEN "1000000",
								
								neighbor64	WHEN "1000001",
								neighbor65	WHEN "1000010",
								neighbor66	WHEN "1000011",
								neighbor67	WHEN "1000100",
								neighbor68	WHEN "1000101",
								neighbor69	WHEN "1000110",
								neighbor70	WHEN "1000111",
								neighbor71	WHEN "1001000",
								neighbor72	WHEN "1001001",
								neighbor73	WHEN "1001010",
								neighbor74	WHEN "1001011",
								neighbor75	WHEN "1001100",
								neighbor76	WHEN "1001101",
								neighbor77	WHEN "1001110",
								neighbor78	WHEN "1001111",
								neighbor79	WHEN "1010000",
								neighbor80	WHEN "1010001",
								neighbor81	WHEN "1010010",
								neighbor82	WHEN "1010011",
								neighbor83	WHEN "1010100",
								neighbor84	WHEN "1010101",
								neighbor85	WHEN "1010110",
								neighbor86	WHEN "1010111",
								neighbor87	WHEN "1011000",
								neighbor88	WHEN "1011001",
								neighbor89	WHEN "1011010",
								neighbor90	WHEN "1011011",
								neighbor91	WHEN OTHERS;
								
	WITH mux_above SELECT
	neighbor_above1	<=	neighbor1	WHEN "0000000",
								neighbor2	WHEN "0000001",
								neighbor3	WHEN "0000010",
								neighbor4	WHEN "0000011",
								neighbor5	WHEN "0000100",
								neighbor6	WHEN "0000101",
								neighbor7	WHEN "0000110",
								neighbor8	WHEN "0000111",
								neighbor9	WHEN "0001000",
								neighbor10	WHEN "0001001",
								neighbor11	WHEN "0001010",
								neighbor12	WHEN "0001011",
								neighbor13	WHEN "0001100",
								neighbor14	WHEN "0001101",
								neighbor15	WHEN "0001110",
								neighbor16	WHEN "0001111",
								neighbor17	WHEN "0010000",
								neighbor18	WHEN "0010001",
								neighbor19	WHEN "0010010",
								neighbor20	WHEN "0010011",
								neighbor21	WHEN "0010100",
								neighbor22	WHEN "0010101",
								neighbor23	WHEN "0010110",
								neighbor24	WHEN "0010111",
								neighbor25	WHEN "0011000",
								neighbor26	WHEN "0011001",
								neighbor27	WHEN "0011010",
								neighbor28	WHEN "0011011",
								neighbor29	WHEN "0011100",
								neighbor30	WHEN "0011101",
								neighbor31	WHEN "0011110",
								neighbor32	WHEN "0011111",
								neighbor33	WHEN "0100000",
								neighbor34	WHEN "0100001",
								neighbor35	WHEN "0100010",
								neighbor36	WHEN "0100011",
								neighbor37	WHEN "0100100",
								neighbor38	WHEN "0100101",
								neighbor39	WHEN "0100110",
								neighbor40	WHEN "0100111",
								neighbor41	WHEN "0101000",
								neighbor42	WHEN "0101001",
								neighbor43	WHEN "0101010",
								neighbor44	WHEN "0101011",
								neighbor45	WHEN "0101100",
								neighbor46	WHEN "0101101",
								neighbor47	WHEN "0101110",
								neighbor48	WHEN "0101111",
								neighbor49	WHEN "0110000",
								neighbor50	WHEN "0110001",
								neighbor51	WHEN "0110010",
								neighbor52	WHEN "0110011",
								neighbor53	WHEN "0110100",
								neighbor54	WHEN "0110101",
								neighbor55	WHEN "0110110",
								neighbor56	WHEN "0110111",
								neighbor57	WHEN "0111000",
								neighbor58	WHEN "0111001",
								neighbor59	WHEN "0111010",
								neighbor60	WHEN "0111011",
								neighbor61	WHEN "0111100",
								neighbor62	WHEN "0111101",
								neighbor63	WHEN "0111110",
								
								neighborDC	WHEN "0111111",
								
								neighbor64	WHEN "1000000",
								neighbor65	WHEN "1000001",
								neighbor66	WHEN "1000010",
								neighbor67	WHEN "1000011",
								neighbor68	WHEN "1000100",
								neighbor69	WHEN "1000101",
								neighbor70	WHEN "1000110",
								neighbor71	WHEN "1000111",
								neighbor72	WHEN "1001000",
								neighbor73	WHEN "1001001",
								neighbor74	WHEN "1001010",
								neighbor75	WHEN "1001011",
								neighbor76	WHEN "1001100",
								neighbor77	WHEN "1001101",
								neighbor78	WHEN "1001110",
								neighbor79	WHEN "1001111",
								neighbor80	WHEN "1010000",
								neighbor81	WHEN "1010001",
								neighbor82	WHEN "1010010",
								neighbor83	WHEN "1010011",
								neighbor84	WHEN "1010100",
								neighbor85	WHEN "1010101",
								neighbor86	WHEN "1010110",
								neighbor87	WHEN "1010111",
								neighbor88	WHEN "1011000",
								neighbor89	WHEN "1011001",
								neighbor90	WHEN "1011010",
								neighbor91	WHEN "1011011",
								neighbor92	WHEN OTHERS;
								
	WITH mux_above SELECT
	neighbor_above2	<= neighbor2	WHEN "0000000",
								neighbor3	WHEN "0000001",
								neighbor4	WHEN "0000010",
								neighbor5	WHEN "0000011",
								neighbor6	WHEN "0000100",
								neighbor7	WHEN "0000101",
								neighbor8	WHEN "0000110",
								neighbor9	WHEN "0000111",
								neighbor10	WHEN "0001000",
								neighbor11	WHEN "0001001",
								neighbor12	WHEN "0001010",
								neighbor13	WHEN "0001011",
								neighbor14	WHEN "0001100",
								neighbor15	WHEN "0001101",
								neighbor16	WHEN "0001110",
								neighbor17	WHEN "0001111",
								neighbor18	WHEN "0010000",
								neighbor19	WHEN "0010001",
								neighbor20	WHEN "0010010",
								neighbor21	WHEN "0010011",
								neighbor22	WHEN "0010100",
								neighbor23	WHEN "0010101",
								neighbor24	WHEN "0010110",
								neighbor25	WHEN "0010111",
								neighbor26	WHEN "0011000",
								neighbor27	WHEN "0011001",
								neighbor28	WHEN "0011010",
								neighbor29	WHEN "0011011",
								neighbor30	WHEN "0011100",
								neighbor31	WHEN "0011101",
								neighbor32	WHEN "0011110",
								neighbor33	WHEN "0011111",
								neighbor34	WHEN "0100000",
								neighbor35	WHEN "0100001",
								neighbor36	WHEN "0100010",
								neighbor37	WHEN "0100011",
								neighbor38	WHEN "0100100",
								neighbor39	WHEN "0100101",
								neighbor40	WHEN "0100110",
								neighbor41	WHEN "0100111",
								neighbor42	WHEN "0101000",
								neighbor43	WHEN "0101001",
								neighbor44	WHEN "0101010",
								neighbor45	WHEN "0101011",
								neighbor46	WHEN "0101100",
								neighbor47	WHEN "0101101",
								neighbor48	WHEN "0101110",
								neighbor49	WHEN "0101111",
								neighbor50	WHEN "0110000",
								neighbor51	WHEN "0110001",
								neighbor52	WHEN "0110010",
								neighbor53	WHEN "0110011",
								neighbor54	WHEN "0110100",
								neighbor55	WHEN "0110101",
								neighbor56	WHEN "0110110",
								neighbor57	WHEN "0110111",
								neighbor58	WHEN "0111000",
								neighbor59	WHEN "0111001",
								neighbor60	WHEN "0111010",
								neighbor61	WHEN "0111011",
								neighbor62	WHEN "0111100",
								neighbor63	WHEN "0111101",
								neighborDC	WHEN "0111110",
								neighbor64	WHEN "0111111",
								neighbor65	WHEN "1000000",
								neighbor66	WHEN "1000001",
								neighbor67	WHEN "1000010",
								neighbor68	WHEN "1000011",
								neighbor69	WHEN "1000100",
								neighbor70	WHEN "1000101",
								neighbor71	WHEN "1000110",
								neighbor72	WHEN "1000111",
								neighbor73	WHEN "1001000",
								neighbor74	WHEN "1001001",
								neighbor75	WHEN "1001010",
								neighbor76	WHEN "1001011",
								neighbor77	WHEN "1001100",
								neighbor78	WHEN "1001101",
								neighbor79	WHEN "1001110",
								neighbor80	WHEN "1001111",
								neighbor81	WHEN "1010000",
								neighbor82	WHEN "1010001",
								neighbor83	WHEN "1010010",
								neighbor84	WHEN "1010011",
								neighbor85	WHEN "1010100",
								neighbor86	WHEN "1010101",
								neighbor87	WHEN "1010110",
								neighbor88	WHEN "1010111",
								neighbor89	WHEN "1011000",
								neighbor90	WHEN "1011001",
								neighbor91	WHEN "1011010",
								neighbor92	WHEN "1011011",
								neighbor93	WHEN OTHERS;
	
	WITH mux_above SELECT
	neighbor_above3	<=	neighbor3	WHEN "0000000",
								neighbor4	WHEN "0000001",
								neighbor5	WHEN "0000010",
								neighbor6	WHEN "0000011",
								neighbor7	WHEN "0000100",
								neighbor8	WHEN "0000101",
								neighbor9	WHEN "0000110",
								neighbor10	WHEN "0000111",
								neighbor11	WHEN "0001000",
								neighbor12	WHEN "0001001",
								neighbor13	WHEN "0001010",
								neighbor14	WHEN "0001011",
								neighbor15	WHEN "0001100",
								neighbor16	WHEN "0001101",
								neighbor17	WHEN "0001110",
								neighbor18	WHEN "0001111",
								neighbor19	WHEN "0010000",
								neighbor20	WHEN "0010001",
								neighbor21	WHEN "0010010",
								neighbor22	WHEN "0010011",
								neighbor23	WHEN "0010100",
								neighbor24	WHEN "0010101",
								neighbor25	WHEN "0010110",
								neighbor26	WHEN "0010111",
								neighbor27	WHEN "0011000",
								neighbor28	WHEN "0011001",
								neighbor29	WHEN "0011010",
								neighbor30	WHEN "0011011",
								neighbor31	WHEN "0011100",
								neighbor32	WHEN "0011101",
								neighbor33	WHEN "0011110",
								neighbor34	WHEN "0011111",
								neighbor35	WHEN "0100000",
								neighbor36	WHEN "0100001",
								neighbor37	WHEN "0100010",
								neighbor38	WHEN "0100011",
								neighbor39	WHEN "0100100",
								neighbor40	WHEN "0100101",
								neighbor41	WHEN "0100110",
								neighbor42	WHEN "0100111",
								neighbor43	WHEN "0101000",
								neighbor44	WHEN "0101001",
								neighbor45	WHEN "0101010",
								neighbor46	WHEN "0101011",
								neighbor47	WHEN "0101100",
								neighbor48	WHEN "0101101",
								neighbor49	WHEN "0101110",
								neighbor50	WHEN "0101111",
								neighbor51	WHEN "0110000",
								neighbor52	WHEN "0110001",
								neighbor53	WHEN "0110010",
								neighbor54	WHEN "0110011",
								neighbor55	WHEN "0110100",
								neighbor56	WHEN "0110101",
								neighbor57	WHEN "0110110",
								neighbor58	WHEN "0110111",
								neighbor59	WHEN "0111000",
								neighbor60	WHEN "0111001",
								neighbor61	WHEN "0111010",
								neighbor62	WHEN "0111011",
								neighbor63	WHEN "0111100",
								
								neighborDC	WHEN "0111101",
								
								neighbor64	WHEN "0111110",
								neighbor65	WHEN "0111111",
								neighbor66	WHEN "1000000",
								neighbor67	WHEN "1000001",
								neighbor68	WHEN "1000010",
								neighbor69	WHEN "1000011",
								neighbor70	WHEN "1000100",
								neighbor71	WHEN "1000101",
								neighbor72	WHEN "1000110",
								neighbor73	WHEN "1000111",
								neighbor74	WHEN "1001000",
								neighbor75	WHEN "1001001",
								neighbor76	WHEN "1001010",
								neighbor77	WHEN "1001011",
								neighbor78	WHEN "1001100",
								neighbor79	WHEN "1001101",
								neighbor80	WHEN "1001110",
								neighbor81	WHEN "1001111",
								neighbor82	WHEN "1010000",
								neighbor83	WHEN "1010001",
								neighbor84	WHEN "1010010",
								neighbor85	WHEN "1010011",
								neighbor86	WHEN "1010100",
								neighbor87	WHEN "1010101",
								neighbor88	WHEN "1010110",
								neighbor89	WHEN "1010111",
								neighbor90	WHEN "1011000",
								neighbor91	WHEN "1011001",
								neighbor92	WHEN "1011010",
								neighbor93	WHEN "1011011",
								neighbor94	WHEN OTHERS;
								
	
	WITH mux_above SELECT
	neighbor_above4	<=	neighbor4	WHEN "0000000",
								neighbor5	WHEN "0000001",
								neighbor6	WHEN "0000010",
								neighbor7	WHEN "0000011",
								neighbor8	WHEN "0000100",
								neighbor9	WHEN "0000101",
								neighbor10	WHEN "0000110",
								neighbor11	WHEN "0000111",
								neighbor12	WHEN "0001000",
								neighbor13	WHEN "0001001",
								neighbor14	WHEN "0001010",
								neighbor15	WHEN "0001011",
								neighbor16	WHEN "0001100",
								neighbor17	WHEN "0001101",
								neighbor18	WHEN "0001110",
								neighbor19	WHEN "0001111",
								neighbor20	WHEN "0010000",
								neighbor21	WHEN "0010001",
								neighbor22	WHEN "0010010",
								neighbor23	WHEN "0010011",
								neighbor24	WHEN "0010100",
								neighbor25	WHEN "0010101",
								neighbor26	WHEN "0010110",
								neighbor27	WHEN "0010111",
								neighbor28	WHEN "0011000",
								neighbor29	WHEN "0011001",
								neighbor30	WHEN "0011010",
								neighbor31	WHEN "0011011",
								neighbor32	WHEN "0011100",
								neighbor33	WHEN "0011101",
								neighbor34	WHEN "0011110",
								neighbor35	WHEN "0011111",
								neighbor36	WHEN "0100000",
								neighbor37	WHEN "0100001",
								neighbor38	WHEN "0100010",
								neighbor39	WHEN "0100011",
								neighbor40	WHEN "0100100",
								neighbor41	WHEN "0100101",
								neighbor42	WHEN "0100110",
								neighbor43	WHEN "0100111",
								neighbor44	WHEN "0101000",
								neighbor45	WHEN "0101001",
								neighbor46	WHEN "0101010",
								neighbor47	WHEN "0101011",
								neighbor48	WHEN "0101100",
								neighbor49	WHEN "0101101",
								neighbor50	WHEN "0101110",
								neighbor51	WHEN "0101111",
								neighbor52	WHEN "0110000",
								neighbor53	WHEN "0110001",
								neighbor54	WHEN "0110010",
								neighbor55	WHEN "0110011",
								neighbor56	WHEN "0110100",
								neighbor57	WHEN "0110101",
								neighbor58	WHEN "0110110",
								neighbor59	WHEN "0110111",
								neighbor60	WHEN "0111000",
								neighbor61	WHEN "0111001",
								neighbor62	WHEN "0111010",
								neighbor63	WHEN "0111011",
								
								neighborDC	WHEN "0111100",
								
								neighbor64	WHEN "0111101",
								neighbor65	WHEN "0111110",
								neighbor66	WHEN "0111111",
								neighbor67	WHEN "1000000",
								neighbor68	WHEN "1000001",
								neighbor69	WHEN "1000010",
								neighbor70	WHEN "1000011",
								neighbor71	WHEN "1000100",
								neighbor72	WHEN "1000101",
								neighbor73	WHEN "1000110",
								neighbor74	WHEN "1000111",
								neighbor75	WHEN "1001000",
								neighbor76	WHEN "1001001",
								neighbor77	WHEN "1001010",
								neighbor78	WHEN "1001011",
								neighbor79	WHEN "1001100",
								neighbor80	WHEN "1001101",
								neighbor81	WHEN "1001110",
								neighbor82	WHEN "1001111",
								neighbor83	WHEN "1010000",
								neighbor84	WHEN "1010001",
								neighbor85	WHEN "1010010",
								neighbor86	WHEN "1010011",
								neighbor87	WHEN "1010100",
								neighbor88	WHEN "1010101",
								neighbor89	WHEN "1010110",
								neighbor90	WHEN "1010111",
								neighbor91	WHEN "1011000",
								neighbor92	WHEN "1011001",
								neighbor93	WHEN "1011010",
								neighbor94	WHEN "1011011",
								neighbor95	WHEN OTHERS;
	
	WITH mux_left SELECT
	neighbor_left0 <=	neighbor32	WHEN "0000000",
							neighbor33	WHEN "0000001",
							neighbor34	WHEN "0000010",
							neighbor35	WHEN "0000011",
							neighbor36	WHEN "0000100",
							neighbor37	WHEN "0000101",
							neighbor38	WHEN "0000110",
							neighbor39	WHEN "0000111",
							neighbor40	WHEN "0001000",
							neighbor41	WHEN "0001001",
							neighbor42	WHEN "0001010",
							neighbor43	WHEN "0001011",
							neighbor44	WHEN "0001100",
							neighbor45	WHEN "0001101",
							neighbor46	WHEN "0001110",
							neighbor47	WHEN "0001111",
							neighbor48	WHEN "0010000",
							neighbor49	WHEN "0010001",
							neighbor50	WHEN "0010010",
							neighbor51	WHEN "0010011",
							neighbor52	WHEN "0010100",
							neighbor53	WHEN "0010101",
							neighbor54	WHEN "0010110",
							neighbor55	WHEN "0010111",
							neighbor56	WHEN "0011000",
							neighbor57	WHEN "0011001",
							neighbor58	WHEN "0011010",
							neighbor59	WHEN "0011011",
							neighbor60	WHEN "0011100",
							neighbor61	WHEN "0011101",
							neighbor62	WHEN "0011110",
							neighbor63	WHEN "0011111",
							
							neighborDC	WHEN "0100000",
							
							neighbor64	WHEN "0100001",
							neighbor65	WHEN "0100010",
							neighbor66	WHEN "0100011",
							neighbor67	WHEN "0100100",
							neighbor68	WHEN "0100101",
							neighbor69	WHEN "0100110",
							neighbor70	WHEN "0100111",
							neighbor71	WHEN "0101000",
							neighbor72	WHEN "0101001",
							neighbor73	WHEN "0101010",
							neighbor74	WHEN "0101011",
							neighbor75	WHEN "0101100",
							neighbor76	WHEN "0101101",
							neighbor77	WHEN "0101110",
							neighbor78	WHEN "0101111",
							neighbor79	WHEN "0110000",
							neighbor80	WHEN "0110001",
							neighbor81	WHEN "0110010",
							neighbor82	WHEN "0110011",
							neighbor83	WHEN "0110100",
							neighbor84	WHEN "0110101",
							neighbor85	WHEN "0110110",
							neighbor86	WHEN "0110111",
							neighbor87	WHEN "0111000",
							neighbor88	WHEN "0111001",
							neighbor89	WHEN "0111010",
							neighbor90	WHEN "0111011",
							neighbor91	WHEN "0111100",
							neighbor92	WHEN "0111101",
							neighbor93	WHEN "0111110",
							neighbor94	WHEN "0111111",
							neighbor95	WHEN "1000000",
							neighbor96	WHEN "1000001",
							neighbor97	WHEN "1000010",
							neighbor98	WHEN "1000011",
							neighbor99	WHEN "1000100",
							neighbor100	WHEN "1000101",
							neighbor101	WHEN "1000110",
							neighbor102	WHEN "1000111",
							neighbor103	WHEN "1001000",
							neighbor104	WHEN "1001001",
							neighbor105	WHEN "1001010",
							neighbor106	WHEN "1001011",
							neighbor107	WHEN "1001100",
							neighbor108	WHEN "1001101",
							neighbor109	WHEN "1001110",
							neighbor110	WHEN "1001111",
							neighbor111	WHEN "1010000",
							neighbor112	WHEN "1010001",
							neighbor113	WHEN "1010010",
							neighbor114	WHEN "1010011",
							neighbor115	WHEN "1010100",
							neighbor116	WHEN "1010101",
							neighbor117	WHEN "1010110",
							neighbor118	WHEN "1010111",
							neighbor119	WHEN "1011000",
							neighbor120	WHEN "1011001",
							neighbor121	WHEN "1011010",
							neighbor122	WHEN "1011011",
							neighbor123	WHEN OTHERS;
							
	WITH mux_left SELECT
	neighbor_left1 <=	neighbor33	WHEN "0000000",
							neighbor34	WHEN "0000001",
							neighbor35	WHEN "0000010",
							neighbor36	WHEN "0000011",
							neighbor37	WHEN "0000100",
							neighbor38	WHEN "0000101",
							neighbor39	WHEN "0000110",
							neighbor40	WHEN "0000111",
							neighbor41	WHEN "0001000",
							neighbor42	WHEN "0001001",
							neighbor43	WHEN "0001010",
							neighbor44	WHEN "0001011",
							neighbor45	WHEN "0001100",
							neighbor46	WHEN "0001101",
							neighbor47	WHEN "0001110",
							neighbor48	WHEN "0001111",
							neighbor49	WHEN "0010000",
							neighbor50	WHEN "0010001",
							neighbor51	WHEN "0010010",
							neighbor52	WHEN "0010011",
							neighbor53	WHEN "0010100",
							neighbor54	WHEN "0010101",
							neighbor55	WHEN "0010110",
							neighbor56	WHEN "0010111",
							neighbor57	WHEN "0011000",
							neighbor58	WHEN "0011001",
							neighbor59	WHEN "0011010",
							neighbor60	WHEN "0011011",
							neighbor61	WHEN "0011100",
							neighbor62	WHEN "0011101",
							neighbor63	WHEN "0011110",
							neighborDC	WHEN "0011111",
							neighbor64	WHEN "0100000",
							neighbor65	WHEN "0100001",
							neighbor66	WHEN "0100010",
							neighbor67	WHEN "0100011",
							neighbor68	WHEN "0100100",
							neighbor69	WHEN "0100101",
							neighbor70	WHEN "0100110",
							neighbor71	WHEN "0100111",
							neighbor72	WHEN "0101000",
							neighbor73	WHEN "0101001",
							neighbor74	WHEN "0101010",
							neighbor75	WHEN "0101011",
							neighbor76	WHEN "0101100",
							neighbor77	WHEN "0101101",
							neighbor78	WHEN "0101110",
							neighbor79	WHEN "0101111",
							neighbor80	WHEN "0110000",
							neighbor81	WHEN "0110001",
							neighbor82	WHEN "0110010",
							neighbor83	WHEN "0110011",
							neighbor84	WHEN "0110100",
							neighbor85	WHEN "0110101",
							neighbor86	WHEN "0110110",
							neighbor87	WHEN "0110111",
							neighbor88	WHEN "0111000",
							neighbor89	WHEN "0111001",
							neighbor90	WHEN "0111010",
							neighbor91	WHEN "0111011",
							neighbor92	WHEN "0111100",
							neighbor93	WHEN "0111101",
							neighbor94	WHEN "0111110",
							neighbor95	WHEN "0111111",
							neighbor96	WHEN "1000000",
							neighbor97	WHEN "1000001",
							neighbor98	WHEN "1000010",
							neighbor99	WHEN "1000011",
							neighbor100	WHEN "1000100",
							neighbor101	WHEN "1000101",
							neighbor102	WHEN "1000110",
							neighbor103	WHEN "1000111",
							neighbor104	WHEN "1001000",
							neighbor105	WHEN "1001001",
							neighbor106	WHEN "1001010",
							neighbor107	WHEN "1001011",
							neighbor108	WHEN "1001100",
							neighbor109	WHEN "1001101",
							neighbor110	WHEN "1001110",
							neighbor111	WHEN "1001111",
							neighbor112	WHEN "1010000",
							neighbor113	WHEN "1010001",
							neighbor114	WHEN "1010010",
							neighbor115	WHEN "1010011",
							neighbor116	WHEN "1010100",
							neighbor117	WHEN "1010101",
							neighbor118	WHEN "1010110",
							neighbor119	WHEN "1010111",
							neighbor120	WHEN "1011000",
							neighbor121	WHEN "1011001",
							neighbor122	WHEN "1011010",
							neighbor123	WHEN "1011011",
							neighbor124	WHEN OTHERS;
	
	WITH mux_left SELECT
	neighbor_left2 <=	neighbor34	WHEN "0000000",
							neighbor35	WHEN "0000001",
							neighbor36	WHEN "0000010",
							neighbor37	WHEN "0000011",
							neighbor38	WHEN "0000100",
							neighbor39	WHEN "0000101",
							neighbor40	WHEN "0000110",
							neighbor41	WHEN "0000111",
							neighbor42	WHEN "0001000",
							neighbor43	WHEN "0001001",
							neighbor44	WHEN "0001010",
							neighbor45	WHEN "0001011",
							neighbor46	WHEN "0001100",
							neighbor47	WHEN "0001101",
							neighbor48	WHEN "0001110",
							neighbor49	WHEN "0001111",
							neighbor50	WHEN "0010000",
							neighbor51	WHEN "0010001",
							neighbor52	WHEN "0010010",
							neighbor53	WHEN "0010011",
							neighbor54	WHEN "0010100",
							neighbor55	WHEN "0010101",
							neighbor56	WHEN "0010110",
							neighbor57	WHEN "0010111",
							neighbor58	WHEN "0011000",
							neighbor59	WHEN "0011001",
							neighbor60	WHEN "0011010",
							neighbor61	WHEN "0011011",
							neighbor62	WHEN "0011100",
							neighbor63	WHEN "0011101",
							neighborDC	WHEN "0011110",
							neighbor64	WHEN "0011111",
							neighbor65	WHEN "0100000",
							neighbor66	WHEN "0100001",
							neighbor67	WHEN "0100010",
							neighbor68	WHEN "0100011",
							neighbor69	WHEN "0100100",
							neighbor70	WHEN "0100101",
							neighbor71	WHEN "0100110",
							neighbor72	WHEN "0100111",
							neighbor73	WHEN "0101000",
							neighbor74	WHEN "0101001",
							neighbor75	WHEN "0101010",
							neighbor76	WHEN "0101011",
							neighbor77	WHEN "0101100",
							neighbor78	WHEN "0101101",
							neighbor79	WHEN "0101110",
							neighbor80	WHEN "0101111",
							neighbor81	WHEN "0110000",
							neighbor82	WHEN "0110001",
							neighbor83	WHEN "0110010",
							neighbor84	WHEN "0110011",
							neighbor85	WHEN "0110100",
							neighbor86	WHEN "0110101",
							neighbor87	WHEN "0110110",
							neighbor88	WHEN "0110111",
							neighbor89	WHEN "0111000",
							neighbor90	WHEN "0111001",
							neighbor91	WHEN "0111010",
							neighbor92	WHEN "0111011",
							neighbor93	WHEN "0111100",
							neighbor94	WHEN "0111101",
							neighbor95	WHEN "0111110",
							neighbor96	WHEN "0111111",
							neighbor97	WHEN "1000000",
							neighbor98	WHEN "1000001",
							neighbor99	WHEN "1000010",
							neighbor100	WHEN "1000011",
							neighbor101	WHEN "1000100",
							neighbor102	WHEN "1000101",
							neighbor103	WHEN "1000110",
							neighbor104	WHEN "1000111",
							neighbor105	WHEN "1001000",
							neighbor106	WHEN "1001001",
							neighbor107	WHEN "1001010",
							neighbor108	WHEN "1001011",
							neighbor109	WHEN "1001100",
							neighbor110	WHEN "1001101",
							neighbor111	WHEN "1001110",
							neighbor112	WHEN "1001111",
							neighbor113	WHEN "1010000",
							neighbor114	WHEN "1010001",
							neighbor115	WHEN "1010010",
							neighbor116	WHEN "1010011",
							neighbor117	WHEN "1010100",
							neighbor118	WHEN "1010101",
							neighbor119	WHEN "1010110",
							neighbor120	WHEN "1010111",
							neighbor121	WHEN "1011000",
							neighbor122	WHEN "1011001",
							neighbor123	WHEN "1011010",
							neighbor124	WHEN "1011011",
							neighbor125	WHEN OTHERS;
							
	WITH mux_left SELECT
	neighbor_left3 <=	neighbor35	WHEN "0000000",
							neighbor36	WHEN "0000001",
							neighbor37	WHEN "0000010",
							neighbor38	WHEN "0000011",
							neighbor39	WHEN "0000100",
							neighbor40	WHEN "0000101",
							neighbor41	WHEN "0000110",
							neighbor42	WHEN "0000111",
							neighbor43	WHEN "0001000",
							neighbor44	WHEN "0001001",
							neighbor45	WHEN "0001010",
							neighbor46	WHEN "0001011",
							neighbor47	WHEN "0001100",
							neighbor48	WHEN "0001101",
							neighbor49	WHEN "0001110",
							neighbor50	WHEN "0001111",
							neighbor51	WHEN "0010000",
							neighbor52	WHEN "0010001",
							neighbor53	WHEN "0010010",
							neighbor54	WHEN "0010011",
							neighbor55	WHEN "0010100",
							neighbor56	WHEN "0010101",
							neighbor57	WHEN "0010110",
							neighbor58	WHEN "0010111",
							neighbor59	WHEN "0011000",
							neighbor60	WHEN "0011001",
							neighbor61	WHEN "0011010",
							neighbor62	WHEN "0011011",
							neighbor63	WHEN "0011100",
							neighborDC	WHEN "0011101",
							neighbor64	WHEN "0011110",
							neighbor65	WHEN "0011111",
							neighbor66	WHEN "0100000",
							neighbor67	WHEN "0100001",
							neighbor68	WHEN "0100010",
							neighbor69	WHEN "0100011",
							neighbor70	WHEN "0100100",
							neighbor71	WHEN "0100101",
							neighbor72	WHEN "0100110",
							neighbor73	WHEN "0100111",
							neighbor74	WHEN "0101000",
							neighbor75	WHEN "0101001",
							neighbor76	WHEN "0101010",
							neighbor77	WHEN "0101011",
							neighbor78	WHEN "0101100",
							neighbor79	WHEN "0101101",
							neighbor80	WHEN "0101110",
							neighbor81	WHEN "0101111",
							neighbor82	WHEN "0110000",
							neighbor83	WHEN "0110001",
							neighbor84	WHEN "0110010",
							neighbor85	WHEN "0110011",
							neighbor86	WHEN "0110100",
							neighbor87	WHEN "0110101",
							neighbor88	WHEN "0110110",
							neighbor89	WHEN "0110111",
							neighbor90	WHEN "0111000",
							neighbor91	WHEN "0111001",
							neighbor92	WHEN "0111010",
							neighbor93	WHEN "0111011",
							neighbor94	WHEN "0111100",
							neighbor95	WHEN "0111101",
							neighbor96	WHEN "0111110",
							neighbor97	WHEN "0111111",
							neighbor98	WHEN "1000000",
							neighbor99	WHEN "1000001",
							neighbor100	WHEN "1000010",
							neighbor101	WHEN "1000011",
							neighbor102	WHEN "1000100",
							neighbor103	WHEN "1000101",
							neighbor104	WHEN "1000110",
							neighbor105	WHEN "1000111",
							neighbor106	WHEN "1001000",
							neighbor107	WHEN "1001001",
							neighbor108	WHEN "1001010",
							neighbor109	WHEN "1001011",
							neighbor110	WHEN "1001100",
							neighbor111	WHEN "1001101",
							neighbor112	WHEN "1001110",
							neighbor113	WHEN "1001111",
							neighbor114	WHEN "1010000",
							neighbor115	WHEN "1010001",
							neighbor116	WHEN "1010010",
							neighbor117	WHEN "1010011",
							neighbor118	WHEN "1010100",
							neighbor119	WHEN "1010101",
							neighbor120	WHEN "1010110",
							neighbor121	WHEN "1010111",
							neighbor122	WHEN "1011000",
							neighbor123	WHEN "1011001",
							neighbor124	WHEN "1011010",
							neighbor125	WHEN "1011011",
							neighbor126	WHEN OTHERS;
	
	WITH mux_left SELECT
	neighbor_left4 <=	neighbor36	WHEN "0000000",
							neighbor37	WHEN "0000001",
							neighbor38	WHEN "0000010",
							neighbor39	WHEN "0000011",
							neighbor40	WHEN "0000100",
							neighbor41	WHEN "0000101",
							neighbor42	WHEN "0000110",
							neighbor43	WHEN "0000111",
							neighbor44	WHEN "0001000",
							neighbor45	WHEN "0001001",
							neighbor46	WHEN "0001010",
							neighbor47	WHEN "0001011",
							neighbor48	WHEN "0001100",
							neighbor49	WHEN "0001101",
							neighbor50	WHEN "0001110",
							neighbor51	WHEN "0001111",
							neighbor52	WHEN "0010000",
							neighbor53	WHEN "0010001",
							neighbor54	WHEN "0010010",
							neighbor55	WHEN "0010011",
							neighbor56	WHEN "0010100",
							neighbor57	WHEN "0010101",
							neighbor58	WHEN "0010110",
							neighbor59	WHEN "0010111",
							neighbor60	WHEN "0011000",
							neighbor61	WHEN "0011001",
							neighbor62	WHEN "0011010",
							neighbor63	WHEN "0011011",
							neighborDC	WHEN "0011100",
							neighbor64	WHEN "0011101",
							neighbor65	WHEN "0011110",
							neighbor66	WHEN "0011111",
							neighbor67	WHEN "0100000",
							neighbor68	WHEN "0100001",
							neighbor69	WHEN "0100010",
							neighbor70	WHEN "0100011",
							neighbor71	WHEN "0100100",
							neighbor72	WHEN "0100101",
							neighbor73	WHEN "0100110",
							neighbor74	WHEN "0100111",
							neighbor75	WHEN "0101000",
							neighbor76	WHEN "0101001",
							neighbor77	WHEN "0101010",
							neighbor78	WHEN "0101011",
							neighbor79	WHEN "0101100",
							neighbor80	WHEN "0101101",
							neighbor81	WHEN "0101110",
							neighbor82	WHEN "0101111",
							neighbor83	WHEN "0110000",
							neighbor84	WHEN "0110001",
							neighbor85	WHEN "0110010",
							neighbor86	WHEN "0110011",
							neighbor87	WHEN "0110100",
							neighbor88	WHEN "0110101",
							neighbor89	WHEN "0110110",
							neighbor90	WHEN "0110111",
							neighbor91	WHEN "0111000",
							neighbor92	WHEN "0111001",
							neighbor93	WHEN "0111010",
							neighbor94	WHEN "0111011",
							neighbor95	WHEN "0111100",
							neighbor96	WHEN "0111101",
							neighbor97	WHEN "0111110",
							neighbor98	WHEN "0111111",
							neighbor99	WHEN "1000000",
							neighbor100	WHEN "1000001",
							neighbor101	WHEN "1000010",
							neighbor102	WHEN "1000011",
							neighbor103	WHEN "1000100",
							neighbor104	WHEN "1000101",
							neighbor105	WHEN "1000110",
							neighbor106	WHEN "1000111",
							neighbor107	WHEN "1001000",
							neighbor108	WHEN "1001001",
							neighbor109	WHEN "1001010",
							neighbor110	WHEN "1001011",
							neighbor111	WHEN "1001100",
							neighbor112	WHEN "1001101",
							neighbor113	WHEN "1001110",
							neighbor114	WHEN "1001111",
							neighbor115	WHEN "1010000",
							neighbor116	WHEN "1010001",
							neighbor117	WHEN "1010010",
							neighbor118	WHEN "1010011",
							neighbor119	WHEN "1010100",
							neighbor120	WHEN "1010101",
							neighbor121	WHEN "1010110",
							neighbor122	WHEN "1010111",
							neighbor123	WHEN "1011000",
							neighbor124	WHEN "1011001",
							neighbor125	WHEN "1011010",
							neighbor126	WHEN "1011011",
							neighbor127	WHEN OTHERS;
							
END behavior;