LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;

ENTITY neighbor_buffer IS
	GENERIC (n: INTEGER:= 8);
	PORT (
		clk,reset		: IN STD_LOGIC;
		enable			: IN STD_LOGIC;
		mux_above		: IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		mux_left			: IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		input_sample	: IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		neighbor_above0: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		neighbor_above1: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		neighbor_above2: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		neighbor_above3: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		neighbor_above4: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		neighbor_left0	: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		neighbor_left1	: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		neighbor_left2	: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		neighbor_left3	: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		neighbor_left4	: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0)
		);
END neighbor_buffer;

ARCHITECTURE behavior OF neighbor_buffer IS

SIGNAL	neighbor0, neighbor1, neighbor2, neighbor3, neighbor4, neighbor5, neighbor6, neighbor7,
			neighbor8, neighbor9, neighbor10,neighbor11,neighbor12,neighbor13,neighbor14,neighbor15,
			neighbor16,neighbor17,neighbor18,neighbor19,neighbor20,neighbor21,neighbor22,neighbor23,
			neighbor24,neighbor25,neighbor26,neighbor27,neighbor28,neighbor29,neighbor30,neighbor31,
			neighbor32,neighbor33,neighbor34,neighbor35,neighbor36,neighbor37,neighbor38,neighbor39,
			neighbor40,neighbor41,neighbor42,neighbor43,neighbor44,neighbor45,neighbor46,neighbor47,
			neighbor48,neighbor49,neighbor50,neighbor51,neighbor52,neighbor53,neighbor54,neighbor55,
			neighbor56,neighbor57,neighbor58,neighbor59,neighbor60,neighbor61,neighbor62,neighbor63,
			neighborDC,
			neighbor64,neighbor65,neighbor66,neighbor67,neighbor68,neighbor69,neighbor70,neighbor71,
			neighbor72,neighbor73,neighbor74,neighbor75,neighbor76,neighbor77,neighbor78,neighbor79,
			neighbor80,neighbor81,neighbor82,neighbor83,neighbor84,neighbor85,neighbor86,neighbor87,
			neighbor88,neighbor89,neighbor90,neighbor91,neighbor92,neighbor93,neighbor94,neighbor95,
			neighbor96, neighbor97, neighbor98, neighbor99, neighbor100,neighbor101,neighbor102,neighbor103,
			neighbor104,neighbor105,neighbor106,neighbor107,neighbor108,neighbor109,neighbor110,neighbor111,
			neighbor112,neighbor113,neighbor114,neighbor115,neighbor116,neighbor117,neighbor118,neighbor119,
			neighbor120,neighbor121,neighbor122,neighbor123,neighbor124,neighbor125,neighbor126,neighbor127
			: STD_LOGIC_VECTOR (n-1 DOWNTO 0);

BEGIN

	PROCESS (clk,reset)
	BEGIN
		IF reset = '1' THEN
			neighbor0 <= (OTHERS=>'0');
			neighbor1 <= (OTHERS=>'0');
			neighbor2 <= (OTHERS=>'0');
			neighbor3 <= (OTHERS=>'0');
			neighbor4 <= (OTHERS=>'0');
			neighbor5 <= (OTHERS=>'0');
			neighbor6 <= (OTHERS=>'0');
			neighbor7 <= (OTHERS=>'0');
			neighbor8 <= (OTHERS=>'0');
			neighbor9 <= (OTHERS=>'0');
			neighbor10 <= (OTHERS=>'0');
			neighbor11 <= (OTHERS=>'0');
			neighbor12 <= (OTHERS=>'0');
			neighbor13 <= (OTHERS=>'0');
			neighbor14 <= (OTHERS=>'0');
			neighbor15 <= (OTHERS=>'0');
			neighbor16 <= (OTHERS=>'0');
			neighbor17 <= (OTHERS=>'0');
			neighbor18 <= (OTHERS=>'0');
			neighbor19 <= (OTHERS=>'0');
			neighbor20 <= (OTHERS=>'0');
			neighbor21 <= (OTHERS=>'0');
			neighbor22 <= (OTHERS=>'0');
			neighbor23 <= (OTHERS=>'0');
			neighbor24 <= (OTHERS=>'0');
			neighbor25 <= (OTHERS=>'0');
			neighbor26 <= (OTHERS=>'0');
			neighbor27 <= (OTHERS=>'0');
			neighbor28 <= (OTHERS=>'0');
			neighbor29 <= (OTHERS=>'0');
			neighbor30 <= (OTHERS=>'0');
			neighbor31 <= (OTHERS=>'0');
			neighbor32 <= (OTHERS=>'0');
			neighbor33 <= (OTHERS=>'0');
			neighbor34 <= (OTHERS=>'0');
			neighbor35 <= (OTHERS=>'0');
			neighbor36 <= (OTHERS=>'0');
			neighbor37 <= (OTHERS=>'0');
			neighbor38 <= (OTHERS=>'0');
			neighbor39 <= (OTHERS=>'0');
			neighbor40 <= (OTHERS=>'0');
			neighbor41 <= (OTHERS=>'0');
			neighbor42 <= (OTHERS=>'0');
			neighbor43 <= (OTHERS=>'0');
			neighbor44 <= (OTHERS=>'0');
			neighbor45 <= (OTHERS=>'0');
			neighbor46 <= (OTHERS=>'0');
			neighbor47 <= (OTHERS=>'0');
			neighbor48 <= (OTHERS=>'0');
			neighbor49 <= (OTHERS=>'0');
			neighbor50 <= (OTHERS=>'0');
			neighbor51 <= (OTHERS=>'0');
			neighbor52 <= (OTHERS=>'0');
			neighbor53 <= (OTHERS=>'0');
			neighbor54 <= (OTHERS=>'0');
			neighbor55 <= (OTHERS=>'0');
			neighbor56 <= (OTHERS=>'0');
			neighbor57 <= (OTHERS=>'0');
			neighbor58 <= (OTHERS=>'0');
			neighbor59 <= (OTHERS=>'0');
			neighbor60 <= (OTHERS=>'0');
			neighbor61 <= (OTHERS=>'0');
			neighbor62 <= (OTHERS=>'0');
			neighbor63 <= (OTHERS=>'0');
			neighborDC <= (OTHERS=>'0');
			neighbor64 <= (OTHERS=>'0');
			neighbor65 <= (OTHERS=>'0');
			neighbor66 <= (OTHERS=>'0');
			neighbor67 <= (OTHERS=>'0');
			neighbor68 <= (OTHERS=>'0');
			neighbor69 <= (OTHERS=>'0');
			neighbor70 <= (OTHERS=>'0');
			neighbor71 <= (OTHERS=>'0');
			neighbor72 <= (OTHERS=>'0');
			neighbor73 <= (OTHERS=>'0');
			neighbor74 <= (OTHERS=>'0');
			neighbor75 <= (OTHERS=>'0');
			neighbor76 <= (OTHERS=>'0');
			neighbor77 <= (OTHERS=>'0');
			neighbor78 <= (OTHERS=>'0');
			neighbor79 <= (OTHERS=>'0');
			neighbor80 <= (OTHERS=>'0');
			neighbor81 <= (OTHERS=>'0');
			neighbor82 <= (OTHERS=>'0');
			neighbor83 <= (OTHERS=>'0');
			neighbor84 <= (OTHERS=>'0');
			neighbor85 <= (OTHERS=>'0');
			neighbor86 <= (OTHERS=>'0');
			neighbor87 <= (OTHERS=>'0');
			neighbor88 <= (OTHERS=>'0');
			neighbor89 <= (OTHERS=>'0');
			neighbor90 <= (OTHERS=>'0');
			neighbor91 <= (OTHERS=>'0');
			neighbor92 <= (OTHERS=>'0');
			neighbor93 <= (OTHERS=>'0');
			neighbor94 <= (OTHERS=>'0');
			neighbor95 <= (OTHERS=>'0');
			neighbor96 <= (OTHERS=>'0');
			neighbor97 <= (OTHERS=>'0');
			neighbor98 <= (OTHERS=>'0');
			neighbor99 <= (OTHERS=>'0');
			neighbor100 <= (OTHERS=>'0');
			neighbor101 <= (OTHERS=>'0');
			neighbor102 <= (OTHERS=>'0');
			neighbor103 <= (OTHERS=>'0');
			neighbor104 <= (OTHERS=>'0');
			neighbor105 <= (OTHERS=>'0');
			neighbor106 <= (OTHERS=>'0');
			neighbor107 <= (OTHERS=>'0');
			neighbor108 <= (OTHERS=>'0');
			neighbor109 <= (OTHERS=>'0');
			neighbor110 <= (OTHERS=>'0');
			neighbor111 <= (OTHERS=>'0');
			neighbor112 <= (OTHERS=>'0');
			neighbor113 <= (OTHERS=>'0');
			neighbor114 <= (OTHERS=>'0');
			neighbor115 <= (OTHERS=>'0');
			neighbor116 <= (OTHERS=>'0');
			neighbor117 <= (OTHERS=>'0');
			neighbor118 <= (OTHERS=>'0');
			neighbor119 <= (OTHERS=>'0');
			neighbor120 <= (OTHERS=>'0');
			neighbor121 <= (OTHERS=>'0');
			neighbor122 <= (OTHERS=>'0');
			neighbor123 <= (OTHERS=>'0');
			neighbor124 <= (OTHERS=>'0');
			neighbor125 <= (OTHERS=>'0');
			neighbor126 <= (OTHERS=>'0');
			neighbor127 <= (OTHERS=>'0');
		ELSIF clk'EVENT AND clk = '1' THEN
			IF enable = '1' THEN
				neighbor0 <= input_sample;
				neighbor1 <= neighbor0;
				neighbor2 <= neighbor1;
				neighbor3 <= neighbor2;
				neighbor4 <= neighbor3;
				neighbor5 <= neighbor4;
				neighbor6 <= neighbor5;
				neighbor7 <= neighbor6;
				neighbor8 <= neighbor7;
				neighbor9 <= neighbor8;
				neighbor10 <= neighbor9;
				neighbor11 <= neighbor10;
				neighbor12 <= neighbor11;
				neighbor13 <= neighbor12;
				neighbor14 <= neighbor13;
				neighbor15 <= neighbor14;
				neighbor16 <= neighbor15;
				neighbor17 <= neighbor16;
				neighbor18 <= neighbor17;
				neighbor19 <= neighbor18;
				neighbor20 <= neighbor19;
				neighbor21 <= neighbor20;
				neighbor22 <= neighbor21;
				neighbor23 <= neighbor22;
				neighbor24 <= neighbor23;
				neighbor25 <= neighbor24;
				neighbor26 <= neighbor25;
				neighbor27 <= neighbor26;
				neighbor28 <= neighbor27;
				neighbor29 <= neighbor28;
				neighbor30 <= neighbor29;
				neighbor31 <= neighbor30;
				neighbor32 <= neighbor31;
				neighbor33 <= neighbor32;
				neighbor34 <= neighbor33;
				neighbor35 <= neighbor34;
				neighbor36 <= neighbor35;
				neighbor37 <= neighbor36;
				neighbor38 <= neighbor37;
				neighbor39 <= neighbor38;
				neighbor40 <= neighbor39;
				neighbor41 <= neighbor40;
				neighbor42 <= neighbor41;
				neighbor43 <= neighbor42;
				neighbor44 <= neighbor43;
				neighbor45 <= neighbor44;
				neighbor46 <= neighbor45;
				neighbor47 <= neighbor46;
				neighbor48 <= neighbor47;
				neighbor49 <= neighbor48;
				neighbor50 <= neighbor49;
				neighbor51 <= neighbor50;
				neighbor52 <= neighbor51;
				neighbor53 <= neighbor52;
				neighbor54 <= neighbor53;
				neighbor55 <= neighbor54;
				neighbor56 <= neighbor55;
				neighbor57 <= neighbor56;
				neighbor58 <= neighbor57;
				neighbor59 <= neighbor58;
				neighbor60 <= neighbor59;
				neighbor61 <= neighbor60;
				neighbor62 <= neighbor61;
				neighbor63 <= neighbor62;
				
				neighborDC <= neighbor63;
				
				neighbor64 <= neighborDC;
				neighbor65 <= neighbor64;
				neighbor66 <= neighbor65;
				neighbor67 <= neighbor66;
				neighbor68 <= neighbor67;
				neighbor69 <= neighbor68;
				neighbor70 <= neighbor69;
				neighbor71 <= neighbor70;
				neighbor72 <= neighbor71;
				neighbor73 <= neighbor72;
				neighbor74 <= neighbor73;
				neighbor75 <= neighbor74;
				neighbor76 <= neighbor75;
				neighbor77 <= neighbor76;
				neighbor78 <= neighbor77;
				neighbor79 <= neighbor78;
				neighbor80 <= neighbor79;
				neighbor81 <= neighbor80;
				neighbor82 <= neighbor81;
				neighbor83 <= neighbor82;
				neighbor84 <= neighbor83;
				neighbor85 <= neighbor84;
				neighbor86 <= neighbor85;
				neighbor87 <= neighbor86;
				neighbor88 <= neighbor87;
				neighbor89 <= neighbor88;
				neighbor90 <= neighbor89;
				neighbor91 <= neighbor90;
				neighbor92 <= neighbor91;
				neighbor93 <= neighbor92;
				neighbor94 <= neighbor93;
				neighbor95 <= neighbor94;
				neighbor96 <= neighbor95;
				neighbor97 <= neighbor96;
				neighbor98 <= neighbor97;
				neighbor99 <= neighbor98;
				neighbor100 <= neighbor99;
				neighbor101 <= neighbor100;
				neighbor102 <= neighbor101;
				neighbor103 <= neighbor102;
				neighbor104 <= neighbor103;
				neighbor105 <= neighbor104;
				neighbor106 <= neighbor105;
				neighbor107 <= neighbor106;
				neighbor108 <= neighbor107;
				neighbor109 <= neighbor108;
				neighbor110 <= neighbor109;
				neighbor111 <= neighbor110;
				neighbor112 <= neighbor111;
				neighbor113 <= neighbor112;
				neighbor114 <= neighbor113;
				neighbor115 <= neighbor114;
				neighbor116 <= neighbor115;
				neighbor117 <= neighbor116;
				neighbor118 <= neighbor117;
				neighbor119 <= neighbor118;
				neighbor120 <= neighbor119;
				neighbor121 <= neighbor120;
				neighbor122 <= neighbor121;
				neighbor123 <= neighbor122;
				neighbor124 <= neighbor123;
				neighbor125 <= neighbor124;
				neighbor126 <= neighbor125;
				neighbor127 <= neighbor126;
			END IF;
		END IF;
	END PROCESS;
	
	WITH mux_above SELECT
	neighbor_above4	<=	neighbor0	WHEN "0000000",
								neighbor0	WHEN "0000001",
								neighbor1	WHEN "0000010",
								neighbor2	WHEN "0000011",
								neighbor3	WHEN "0000100",
								neighbor4	WHEN "0000101",
								neighbor5	WHEN "0000110",
								neighbor6	WHEN "0000111",
								neighbor7	WHEN "0001000",
								neighbor8	WHEN "0001001",
								neighbor9	WHEN "0001010",
								neighbor10	WHEN "0001011",
								neighbor11	WHEN "0001100",
								neighbor12	WHEN "0001101",
								neighbor13	WHEN "0001110",
								neighbor14	WHEN "0001111",
								neighbor15	WHEN "0010000",
								neighbor16	WHEN "0010001",
								neighbor17	WHEN "0010010",
								neighbor18	WHEN "0010011",
								neighbor19	WHEN "0010100",
								neighbor20	WHEN "0010101",
								neighbor21	WHEN "0010110",
								neighbor22	WHEN "0010111",
								neighbor23	WHEN "0011000",
								neighbor24	WHEN "0011001",
								neighbor25	WHEN "0011010",
								neighbor26	WHEN "0011011",
								neighbor27	WHEN "0011100",
								neighbor28	WHEN "0011101",
								neighbor29	WHEN "0011110",
								neighbor30	WHEN "0011111",
								neighbor31	WHEN "0100000",
								neighbor32	WHEN "0100001",
								neighbor33	WHEN "0100010",
								neighbor34	WHEN "0100011",
								neighbor35	WHEN "0100100",
								neighbor36	WHEN "0100101",
								neighbor37	WHEN "0100110",
								neighbor38	WHEN "0100111",
								neighbor39	WHEN "0101000",
								neighbor40	WHEN "0101001",
								neighbor41	WHEN "0101010",
								neighbor42	WHEN "0101011",
								neighbor43	WHEN "0101100",
								neighbor44	WHEN "0101101",
								neighbor45	WHEN "0101110",
								neighbor46	WHEN "0101111",
								neighbor47	WHEN "0110000",
								neighbor48	WHEN "0110001",
								neighbor49	WHEN "0110010",
								neighbor50	WHEN "0110011",
								neighbor51	WHEN "0110100",
								neighbor52	WHEN "0110101",
								neighbor53	WHEN "0110110",
								neighbor54	WHEN "0110111",
								neighbor55	WHEN "0111000",
								neighbor56	WHEN "0111001",
								neighbor57	WHEN "0111010",
								neighbor58	WHEN "0111011",
								neighbor59	WHEN "0111100",
								neighbor60	WHEN "0111101",
								neighbor61	WHEN "0111110",
								neighbor62	WHEN "0111111",
								neighbor63	WHEN "1000000",
								neighborDC	WHEN "1000001",
								neighbor64	WHEN "1000010",
								neighbor65	WHEN "1000011",
								neighbor66	WHEN "1000100",
								neighbor67	WHEN "1000101",
								neighbor68	WHEN "1000110",
								neighbor69	WHEN "1000111",
								neighbor70	WHEN "1001000",
								neighbor71	WHEN "1001001",
								neighbor72	WHEN "1001010",
								neighbor73	WHEN "1001011",
								neighbor74	WHEN "1001100",
								neighbor75	WHEN "1001101",
								neighbor76	WHEN "1001110",
								neighbor77	WHEN "1001111",
								neighbor78	WHEN "1010000",
								neighbor79	WHEN "1010001",
								neighbor80	WHEN "1010010",
								neighbor81	WHEN "1010011",
								neighbor82	WHEN "1010100",
								neighbor83	WHEN "1010101",
								neighbor84	WHEN "1010110",
								neighbor85	WHEN "1010111",
								neighbor86	WHEN "1011000",
								neighbor87	WHEN "1011001",
								neighbor88	WHEN "1011010",
								neighbor89	WHEN "1011011",
								neighbor90	WHEN "1011100",
								neighbor91	WHEN OTHERS;
								
	WITH mux_above SELECT
	neighbor_above3	<=	neighbor0	WHEN "0000000",
								neighbor1	WHEN "0000001",
								neighbor2	WHEN "0000010",
								neighbor3	WHEN "0000011",
								neighbor4	WHEN "0000100",
								neighbor5	WHEN "0000101",
								neighbor6	WHEN "0000110",
								neighbor7	WHEN "0000111",
								neighbor8	WHEN "0001000",
								neighbor9	WHEN "0001001",
								neighbor10	WHEN "0001010",
								neighbor11	WHEN "0001011",
								neighbor12	WHEN "0001100",
								neighbor13	WHEN "0001101",
								neighbor14	WHEN "0001110",
								neighbor15	WHEN "0001111",
								neighbor16	WHEN "0010000",
								neighbor17	WHEN "0010001",
								neighbor18	WHEN "0010010",
								neighbor19	WHEN "0010011",
								neighbor20	WHEN "0010100",
								neighbor21	WHEN "0010101",
								neighbor22	WHEN "0010110",
								neighbor23	WHEN "0010111",
								neighbor24	WHEN "0011000",
								neighbor25	WHEN "0011001",
								neighbor26	WHEN "0011010",
								neighbor27	WHEN "0011011",
								neighbor28	WHEN "0011100",
								neighbor29	WHEN "0011101",
								neighbor30	WHEN "0011110",
								neighbor31	WHEN "0011111",
								neighbor32	WHEN "0100000",
								neighbor33	WHEN "0100001",
								neighbor34	WHEN "0100010",
								neighbor35	WHEN "0100011",
								neighbor36	WHEN "0100100",
								neighbor37	WHEN "0100101",
								neighbor38	WHEN "0100110",
								neighbor39	WHEN "0100111",
								neighbor40	WHEN "0101000",
								neighbor41	WHEN "0101001",
								neighbor42	WHEN "0101010",
								neighbor43	WHEN "0101011",
								neighbor44	WHEN "0101100",
								neighbor45	WHEN "0101101",
								neighbor46	WHEN "0101110",
								neighbor47	WHEN "0101111",
								neighbor48	WHEN "0110000",
								neighbor49	WHEN "0110001",
								neighbor50	WHEN "0110010",
								neighbor51	WHEN "0110011",
								neighbor52	WHEN "0110100",
								neighbor53	WHEN "0110101",
								neighbor54	WHEN "0110110",
								neighbor55	WHEN "0110111",
								neighbor56	WHEN "0111000",
								neighbor57	WHEN "0111001",
								neighbor58	WHEN "0111010",
								neighbor59	WHEN "0111011",
								neighbor60	WHEN "0111100",
								neighbor61	WHEN "0111101",
								neighbor62	WHEN "0111110",
								neighbor63	WHEN "0111111",
								neighborDC	WHEN "1000000",
								neighbor64	WHEN "1000001",
								neighbor65	WHEN "1000010",
								neighbor66	WHEN "1000011",
								neighbor67	WHEN "1000100",
								neighbor68	WHEN "1000101",
								neighbor69	WHEN "1000110",
								neighbor70	WHEN "1000111",
								neighbor71	WHEN "1001000",
								neighbor72	WHEN "1001001",
								neighbor73	WHEN "1001010",
								neighbor74	WHEN "1001011",
								neighbor75	WHEN "1001100",
								neighbor76	WHEN "1001101",
								neighbor77	WHEN "1001110",
								neighbor78	WHEN "1001111",
								neighbor79	WHEN "1010000",
								neighbor80	WHEN "1010001",
								neighbor81	WHEN "1010010",
								neighbor82	WHEN "1010011",
								neighbor83	WHEN "1010100",
								neighbor84	WHEN "1010101",
								neighbor85	WHEN "1010110",
								neighbor86	WHEN "1010111",
								neighbor87	WHEN "1011000",
								neighbor88	WHEN "1011001",
								neighbor89	WHEN "1011010",
								neighbor90	WHEN "1011011",
								neighbor91	WHEN "1011100",
								neighbor92	WHEN OTHERS;
								
	WITH mux_above SELECT
	neighbor_above2	<= neighbor1	WHEN "0000000",
								neighbor2	WHEN "0000001",
								neighbor3	WHEN "0000010",
								neighbor4	WHEN "0000011",
								neighbor5	WHEN "0000100",
								neighbor6	WHEN "0000101",
								neighbor7	WHEN "0000110",
								neighbor8	WHEN "0000111",
								neighbor9	WHEN "0001000",
								neighbor10	WHEN "0001001",
								neighbor11	WHEN "0001010",
								neighbor12	WHEN "0001011",
								neighbor13	WHEN "0001100",
								neighbor14	WHEN "0001101",
								neighbor15	WHEN "0001110",
								neighbor16	WHEN "0001111",
								neighbor17	WHEN "0010000",
								neighbor18	WHEN "0010001",
								neighbor19	WHEN "0010010",
								neighbor20	WHEN "0010011",
								neighbor21	WHEN "0010100",
								neighbor22	WHEN "0010101",
								neighbor23	WHEN "0010110",
								neighbor24	WHEN "0010111",
								neighbor25	WHEN "0011000",
								neighbor26	WHEN "0011001",
								neighbor27	WHEN "0011010",
								neighbor28	WHEN "0011011",
								neighbor29	WHEN "0011100",
								neighbor30	WHEN "0011101",
								neighbor31	WHEN "0011110",
								neighbor32	WHEN "0011111",
								neighbor33	WHEN "0100000",
								neighbor34	WHEN "0100001",
								neighbor35	WHEN "0100010",
								neighbor36	WHEN "0100011",
								neighbor37	WHEN "0100100",
								neighbor38	WHEN "0100101",
								neighbor39	WHEN "0100110",
								neighbor40	WHEN "0100111",
								neighbor41	WHEN "0101000",
								neighbor42	WHEN "0101001",
								neighbor43	WHEN "0101010",
								neighbor44	WHEN "0101011",
								neighbor45	WHEN "0101100",
								neighbor46	WHEN "0101101",
								neighbor47	WHEN "0101110",
								neighbor48	WHEN "0101111",
								neighbor49	WHEN "0110000",
								neighbor50	WHEN "0110001",
								neighbor51	WHEN "0110010",
								neighbor52	WHEN "0110011",
								neighbor53	WHEN "0110100",
								neighbor54	WHEN "0110101",
								neighbor55	WHEN "0110110",
								neighbor56	WHEN "0110111",
								neighbor57	WHEN "0111000",
								neighbor58	WHEN "0111001",
								neighbor59	WHEN "0111010",
								neighbor60	WHEN "0111011",
								neighbor61	WHEN "0111100",
								neighbor62	WHEN "0111101",
								neighbor63	WHEN "0111110",
								neighborDC	WHEN "0111111",
								neighbor64	WHEN "1000000",
								neighbor65	WHEN "1000001",
								neighbor66	WHEN "1000010",
								neighbor67	WHEN "1000011",
								neighbor68	WHEN "1000100",
								neighbor69	WHEN "1000101",
								neighbor70	WHEN "1000110",
								neighbor71	WHEN "1000111",
								neighbor72	WHEN "1001000",
								neighbor73	WHEN "1001001",
								neighbor74	WHEN "1001010",
								neighbor75	WHEN "1001011",
								neighbor76	WHEN "1001100",
								neighbor77	WHEN "1001101",
								neighbor78	WHEN "1001110",
								neighbor79	WHEN "1001111",
								neighbor80	WHEN "1010000",
								neighbor81	WHEN "1010001",
								neighbor82	WHEN "1010010",
								neighbor83	WHEN "1010011",
								neighbor84	WHEN "1010100",
								neighbor85	WHEN "1010101",
								neighbor86	WHEN "1010110",
								neighbor87	WHEN "1010111",
								neighbor88	WHEN "1011000",
								neighbor89	WHEN "1011001",
								neighbor90	WHEN "1011010",
								neighbor91	WHEN "1011011",
								neighbor92	WHEN "1011100",
								neighbor93	WHEN OTHERS;
	
	WITH mux_above SELECT
	neighbor_above1	<=	neighbor2	WHEN "0000000",
								neighbor3	WHEN "0000001",
								neighbor4	WHEN "0000010",
								neighbor5	WHEN "0000011",
								neighbor6	WHEN "0000100",
								neighbor7	WHEN "0000101",
								neighbor8	WHEN "0000110",
								neighbor9	WHEN "0000111",
								neighbor10	WHEN "0001000",
								neighbor11	WHEN "0001001",
								neighbor12	WHEN "0001010",
								neighbor13	WHEN "0001011",
								neighbor14	WHEN "0001100",
								neighbor15	WHEN "0001101",
								neighbor16	WHEN "0001110",
								neighbor17	WHEN "0001111",
								neighbor18	WHEN "0010000",
								neighbor19	WHEN "0010001",
								neighbor20	WHEN "0010010",
								neighbor21	WHEN "0010011",
								neighbor22	WHEN "0010100",
								neighbor23	WHEN "0010101",
								neighbor24	WHEN "0010110",
								neighbor25	WHEN "0010111",
								neighbor26	WHEN "0011000",
								neighbor27	WHEN "0011001",
								neighbor28	WHEN "0011010",
								neighbor29	WHEN "0011011",
								neighbor30	WHEN "0011100",
								neighbor31	WHEN "0011101",
								neighbor32	WHEN "0011110",
								neighbor33	WHEN "0011111",
								neighbor34	WHEN "0100000",
								neighbor35	WHEN "0100001",
								neighbor36	WHEN "0100010",
								neighbor37	WHEN "0100011",
								neighbor38	WHEN "0100100",
								neighbor39	WHEN "0100101",
								neighbor40	WHEN "0100110",
								neighbor41	WHEN "0100111",
								neighbor42	WHEN "0101000",
								neighbor43	WHEN "0101001",
								neighbor44	WHEN "0101010",
								neighbor45	WHEN "0101011",
								neighbor46	WHEN "0101100",
								neighbor47	WHEN "0101101",
								neighbor48	WHEN "0101110",
								neighbor49	WHEN "0101111",
								neighbor50	WHEN "0110000",
								neighbor51	WHEN "0110001",
								neighbor52	WHEN "0110010",
								neighbor53	WHEN "0110011",
								neighbor54	WHEN "0110100",
								neighbor55	WHEN "0110101",
								neighbor56	WHEN "0110110",
								neighbor57	WHEN "0110111",
								neighbor58	WHEN "0111000",
								neighbor59	WHEN "0111001",
								neighbor60	WHEN "0111010",
								neighbor61	WHEN "0111011",
								neighbor62	WHEN "0111100",
								neighbor63	WHEN "0111101",
								neighborDC	WHEN "0111110",
								neighbor64	WHEN "0111111",
								neighbor65	WHEN "1000000",
								neighbor66	WHEN "1000001",
								neighbor67	WHEN "1000010",
								neighbor68	WHEN "1000011",
								neighbor69	WHEN "1000100",
								neighbor70	WHEN "1000101",
								neighbor71	WHEN "1000110",
								neighbor72	WHEN "1000111",
								neighbor73	WHEN "1001000",
								neighbor74	WHEN "1001001",
								neighbor75	WHEN "1001010",
								neighbor76	WHEN "1001011",
								neighbor77	WHEN "1001100",
								neighbor78	WHEN "1001101",
								neighbor79	WHEN "1001110",
								neighbor80	WHEN "1001111",
								neighbor81	WHEN "1010000",
								neighbor82	WHEN "1010001",
								neighbor83	WHEN "1010010",
								neighbor84	WHEN "1010011",
								neighbor85	WHEN "1010100",
								neighbor86	WHEN "1010101",
								neighbor87	WHEN "1010110",
								neighbor88	WHEN "1010111",
								neighbor89	WHEN "1011000",
								neighbor90	WHEN "1011001",
								neighbor91	WHEN "1011010",
								neighbor92	WHEN "1011011",
								neighbor93	WHEN "1011100",
								neighbor94	WHEN OTHERS;
								
	--CABECA!!!!!!
	WITH mux_above SELECT
	neighbor_above0	<=	neighbor3	WHEN "0000000",
								neighbor4	WHEN "0000001",
								neighbor5	WHEN "0000010",
								neighbor6	WHEN "0000011",
								neighbor7	WHEN "0000100",
								neighbor8	WHEN "0000101",
								neighbor9	WHEN "0000110",
								neighbor10	WHEN "0000111",
								neighbor11	WHEN "0001000",
								neighbor12	WHEN "0001001",
								neighbor13	WHEN "0001010",
								neighbor14	WHEN "0001011",
								neighbor15	WHEN "0001100",
								neighbor16	WHEN "0001101",
								neighbor17	WHEN "0001110",
								neighbor18	WHEN "0001111",
								neighbor19	WHEN "0010000",
								neighbor20	WHEN "0010001",
								neighbor21	WHEN "0010010",
								neighbor22	WHEN "0010011",
								neighbor23	WHEN "0010100",
								neighbor24	WHEN "0010101",
								neighbor25	WHEN "0010110",
								neighbor26	WHEN "0010111",
								neighbor27	WHEN "0011000",
								neighbor28	WHEN "0011001",
								neighbor29	WHEN "0011010",
								neighbor30	WHEN "0011011",
								neighbor31	WHEN "0011100",
								neighbor32	WHEN "0011101",
								neighbor33	WHEN "0011110",
								neighbor34	WHEN "0011111",
								neighbor35	WHEN "0100000",
								neighbor36	WHEN "0100001",
								neighbor37	WHEN "0100010",
								neighbor38	WHEN "0100011",
								neighbor39	WHEN "0100100",
								neighbor40	WHEN "0100101",
								neighbor41	WHEN "0100110",
								neighbor42	WHEN "0100111",
								neighbor43	WHEN "0101000",
								neighbor44	WHEN "0101001",
								neighbor45	WHEN "0101010",
								neighbor46	WHEN "0101011",
								neighbor47	WHEN "0101100",
								neighbor48	WHEN "0101101",
								neighbor49	WHEN "0101110",
								neighbor50	WHEN "0101111",
								neighbor51	WHEN "0110000",
								neighbor52	WHEN "0110001",
								neighbor53	WHEN "0110010",
								neighbor54	WHEN "0110011",
								neighbor55	WHEN "0110100",
								neighbor56	WHEN "0110101",
								neighbor57	WHEN "0110110",
								neighbor58	WHEN "0110111",
								neighbor59	WHEN "0111000",
								neighbor60	WHEN "0111001",
								neighbor61	WHEN "0111010",
								neighbor62	WHEN "0111011", --59
								neighbor63	WHEN "0111100", --60
								neighborDC	WHEN "0111101", --61
								neighbor64	WHEN "0111110", --62
								neighbor65	WHEN "0111111",
								neighbor66	WHEN "1000000",
								neighbor67	WHEN "1000001",
								neighbor68	WHEN "1000010",
								neighbor69	WHEN "1000011",
								neighbor70	WHEN "1000100",
								neighbor71	WHEN "1000101",
								neighbor72	WHEN "1000110",
								neighbor73	WHEN "1000111",
								neighbor74	WHEN "1001000",
								neighbor75	WHEN "1001001",
								neighbor76	WHEN "1001010",
								neighbor77	WHEN "1001011",
								neighbor78	WHEN "1001100",
								neighbor79	WHEN "1001101",
								neighbor80	WHEN "1001110",
								neighbor81	WHEN "1001111",
								neighbor82	WHEN "1010000",
								neighbor83	WHEN "1010001",
								neighbor84	WHEN "1010010",
								neighbor85	WHEN "1010011",
								neighbor86	WHEN "1010100",
								neighbor87	WHEN "1010101",
								neighbor88	WHEN "1010110",
								neighbor89	WHEN "1010111",
								neighbor90	WHEN "1011000",
								neighbor91	WHEN "1011001",
								neighbor92	WHEN "1011010",
								neighbor93	WHEN "1011011",
								neighbor94	WHEN "1011100",
								neighbor95	WHEN OTHERS;
	
	WITH mux_left SELECT
	neighbor_left4 <=	neighbor124	WHEN "0000000",
							neighbor123	WHEN "0000001",
							neighbor122	WHEN "0000010",
							neighbor121	WHEN "0000011",
							neighbor120	WHEN "0000100",
							neighbor119	WHEN "0000101",
							neighbor118	WHEN "0000110",
							neighbor117	WHEN "0000111",
							neighbor116	WHEN "0001000",
							neighbor115	WHEN "0001001",
							neighbor114	WHEN "0001010",
							neighbor113	WHEN "0001011",
							neighbor112	WHEN "0001100",
							neighbor111	WHEN "0001101",
							neighbor110	WHEN "0001110",
							neighbor109	WHEN "0001111",
							neighbor108	WHEN "0010000",
							neighbor107	WHEN "0010001",
							neighbor106	WHEN "0010010",
							neighbor105	WHEN "0010011",
							neighbor104	WHEN "0010100",
							neighbor103	WHEN "0010101",
							neighbor102	WHEN "0010110",
							neighbor101	WHEN "0010111",
							neighbor100	WHEN "0011000",
							neighbor99	WHEN "0011001",
							neighbor98	WHEN "0011010",
							neighbor97	WHEN "0011011",
							neighbor96	WHEN "0011100",
							neighbor95	WHEN "0011101",
							neighbor94	WHEN "0011110",
							neighbor93	WHEN "0011111",
							neighbor92	WHEN "0100000",
							neighbor91	WHEN "0100001",
							neighbor90	WHEN "0100010",
							neighbor89	WHEN "0100011",
							neighbor88	WHEN "0100100",
							neighbor87	WHEN "0100101",
							neighbor86	WHEN "0100110",
							neighbor85	WHEN "0100111",
							neighbor84	WHEN "0101000",
							neighbor83	WHEN "0101001",
							neighbor82	WHEN "0101010",
							neighbor81	WHEN "0101011",
							neighbor80	WHEN "0101100",
							neighbor79	WHEN "0101101",
							neighbor78	WHEN "0101110",
							neighbor77	WHEN "0101111",
							neighbor76	WHEN "0110000",
							neighbor75	WHEN "0110001",
							neighbor74	WHEN "0110010",
							neighbor73	WHEN "0110011",
							neighbor72	WHEN "0110100",
							neighbor71	WHEN "0110101",
							neighbor70	WHEN "0110110",
							neighbor69	WHEN "0110111",
							neighbor68	WHEN "0111000",
							neighbor67	WHEN "0111001",
							neighbor66	WHEN "0111010",
							neighbor65	WHEN "0111011",
							neighborDC	WHEN "0111100",
							neighbor64	WHEN "0111101",
							neighbor63	WHEN "0111110",
							neighbor62	WHEN "0111111",
							neighbor61	WHEN "1000000",
							neighbor60	WHEN "1000001",
							neighbor59	WHEN "1000010",
							neighbor58	WHEN "1000011",
							neighbor57	WHEN "1000100",
							neighbor56	WHEN "1000101",
							neighbor55	WHEN "1000110",
							neighbor54	WHEN "1000111",
							neighbor53	WHEN "1001000",
							neighbor52	WHEN "1001001",
							neighbor51	WHEN "1001010",
							neighbor50	WHEN "1001011",
							neighbor49	WHEN "1001100",
							neighbor48	WHEN "1001101",
							neighbor47	WHEN "1001110",
							neighbor46	WHEN "1001111",
							neighbor45	WHEN "1010000",
							neighbor44	WHEN "1010001",
							neighbor43	WHEN "1010010",
							neighbor42	WHEN "1010011",
							neighbor41	WHEN "1010100",
							neighbor40	WHEN "1010101",
							neighbor39	WHEN "1010110",
							neighbor38	WHEN "1010111",
							neighbor37	WHEN "1011000",
							neighbor36	WHEN "1011001",
							neighbor35	WHEN "1011010",
							neighbor34	WHEN "1011011",
							neighbor33	WHEN "1011100",
							neighbor32	WHEN OTHERS;
							
	WITH mux_left SELECT
	neighbor_left3 <=	neighbor125	WHEN "0000000",
							neighbor124	WHEN "0000001",
							neighbor123	WHEN "0000010",
							neighbor122	WHEN "0000011",
							neighbor121	WHEN "0000100",
							neighbor120	WHEN "0000101",
							neighbor119	WHEN "0000110",
							neighbor118	WHEN "0000111",
							neighbor117	WHEN "0001000",
							neighbor116	WHEN "0001001",
							neighbor115	WHEN "0001010",
							neighbor114	WHEN "0001011",
							neighbor113	WHEN "0001100",
							neighbor112	WHEN "0001101",
							neighbor111	WHEN "0001110",
							neighbor110	WHEN "0001111",
							neighbor109	WHEN "0010000",
							neighbor108	WHEN "0010001",
							neighbor107	WHEN "0010010",
							neighbor106	WHEN "0010011",
							neighbor105	WHEN "0010100",
							neighbor104	WHEN "0010101",
							neighbor103	WHEN "0010110",
							neighbor102	WHEN "0010111",
							neighbor101	WHEN "0011000",
							neighbor100	WHEN "0011001",
							neighbor99	WHEN "0011010",
							neighbor98	WHEN "0011011",
							neighbor97	WHEN "0011100",
							neighbor96	WHEN "0011101",
							neighbor95	WHEN "0011110",
							neighbor94	WHEN "0011111",
							neighbor93	WHEN "0100000",
							neighbor92	WHEN "0100001",
							neighbor91	WHEN "0100010",
							neighbor90	WHEN "0100011",
							neighbor89	WHEN "0100100",
							neighbor88	WHEN "0100101",
							neighbor87	WHEN "0100110",
							neighbor86	WHEN "0100111",
							neighbor85	WHEN "0101000",
							neighbor84	WHEN "0101001",
							neighbor83	WHEN "0101010",
							neighbor82	WHEN "0101011",
							neighbor81	WHEN "0101100",
							neighbor80	WHEN "0101101",
							neighbor79	WHEN "0101110",
							neighbor78	WHEN "0101111",
							neighbor77	WHEN "0110000",
							neighbor76	WHEN "0110001",
							neighbor75	WHEN "0110010",
							neighbor74	WHEN "0110011",
							neighbor73	WHEN "0110100",
							neighbor72	WHEN "0110101",
							neighbor71	WHEN "0110110",
							neighbor70	WHEN "0110111",
							neighbor69	WHEN "0111000",
							neighbor68	WHEN "0111001",
							neighbor67	WHEN "0111010",
							neighbor66	WHEN "0111011",
							neighbor65	WHEN "0111100",
							neighborDC	WHEN "0111101",
							neighbor64	WHEN "0111110",
							neighbor63	WHEN "0111111",
							neighbor62	WHEN "1000000",
							neighbor61	WHEN "1000001",
							neighbor60	WHEN "1000010",
							neighbor59	WHEN "1000011",
							neighbor58	WHEN "1000100",
							neighbor57	WHEN "1000101",
							neighbor56	WHEN "1000110",
							neighbor55	WHEN "1000111",
							neighbor54	WHEN "1001000",
							neighbor53	WHEN "1001001",
							neighbor52	WHEN "1001010",
							neighbor51	WHEN "1001011",
							neighbor50	WHEN "1001100",
							neighbor49	WHEN "1001101",
							neighbor48	WHEN "1001110",
							neighbor47	WHEN "1001111",
							neighbor46	WHEN "1010000",
							neighbor45	WHEN "1010001",
							neighbor44	WHEN "1010010",
							neighbor43	WHEN "1010011",
							neighbor42	WHEN "1010100",
							neighbor41	WHEN "1010101",
							neighbor40	WHEN "1010110",
							neighbor39	WHEN "1010111",
							neighbor38	WHEN "1011000",
							neighbor37	WHEN "1011001",
							neighbor36	WHEN "1011010",
							neighbor35	WHEN "1011011",
							neighbor34	WHEN "1011100",
							neighbor33	WHEN OTHERS;
	
	WITH mux_left SELECT
	neighbor_left2 <=	neighbor126	WHEN "0000000",
							neighbor125	WHEN "0000001",
							neighbor124	WHEN "0000010",
							neighbor123	WHEN "0000011",
							neighbor122	WHEN "0000100",
							neighbor121	WHEN "0000101",
							neighbor120	WHEN "0000110",
							neighbor119	WHEN "0000111",
							neighbor118	WHEN "0001000",
							neighbor117	WHEN "0001001",
							neighbor116	WHEN "0001010",
							neighbor115	WHEN "0001011",
							neighbor114	WHEN "0001100",
							neighbor113	WHEN "0001101",
							neighbor112	WHEN "0001110",
							neighbor111	WHEN "0001111",
							neighbor110	WHEN "0010000",
							neighbor109	WHEN "0010001",
							neighbor108	WHEN "0010010",
							neighbor107	WHEN "0010011",
							neighbor106	WHEN "0010100",
							neighbor105	WHEN "0010101",
							neighbor104	WHEN "0010110",
							neighbor103	WHEN "0010111",
							neighbor102	WHEN "0011000",
							neighbor101	WHEN "0011001",
							neighbor100	WHEN "0011010",
							neighbor99	WHEN "0011011",
							neighbor98	WHEN "0011100",
							neighbor97	WHEN "0011101",
							neighbor96	WHEN "0011110",
							neighbor95	WHEN "0011111",
							neighbor94	WHEN "0100000",
							neighbor93	WHEN "0100001",
							neighbor92	WHEN "0100010",
							neighbor91	WHEN "0100011",
							neighbor90	WHEN "0100100",
							neighbor89	WHEN "0100101",
							neighbor88	WHEN "0100110",
							neighbor87	WHEN "0100111",
							neighbor86	WHEN "0101000",
							neighbor85	WHEN "0101001",
							neighbor84	WHEN "0101010",
							neighbor83	WHEN "0101011",
							neighbor82	WHEN "0101100",
							neighbor81	WHEN "0101101",
							neighbor80	WHEN "0101110",
							neighbor79	WHEN "0101111",
							neighbor78	WHEN "0110000",
							neighbor77	WHEN "0110001",
							neighbor76	WHEN "0110010",
							neighbor75	WHEN "0110011",
							neighbor74	WHEN "0110100",
							neighbor73	WHEN "0110101",
							neighbor72	WHEN "0110110",
							neighbor71	WHEN "0110111",
							neighbor70	WHEN "0111000",
							neighbor69	WHEN "0111001",
							neighbor68	WHEN "0111010",
							neighbor67	WHEN "0111011",
							neighbor66	WHEN "0111100",
							neighbor65	WHEN "0111101",
							neighborDC	WHEN "0111110",
							neighbor64	WHEN "0111111",
							neighbor63	WHEN "1000000",
							neighbor62	WHEN "1000001",
							neighbor61	WHEN "1000010",
							neighbor60	WHEN "1000011",
							neighbor59	WHEN "1000100",
							neighbor58	WHEN "1000101",
							neighbor57	WHEN "1000110",
							neighbor56	WHEN "1000111",
							neighbor55	WHEN "1001000",
							neighbor54	WHEN "1001001",
							neighbor53	WHEN "1001010",
							neighbor52	WHEN "1001011",
							neighbor51	WHEN "1001100",
							neighbor50	WHEN "1001101",
							neighbor49	WHEN "1001110",
							neighbor48	WHEN "1001111",
							neighbor47	WHEN "1010000",
							neighbor46	WHEN "1010001",
							neighbor45	WHEN "1010010",
							neighbor44	WHEN "1010011",
							neighbor43	WHEN "1010100",
							neighbor42	WHEN "1010101",
							neighbor41	WHEN "1010110",
							neighbor40	WHEN "1010111",
							neighbor39	WHEN "1011000",
							neighbor38	WHEN "1011001",
							neighbor37	WHEN "1011010",
							neighbor36	WHEN "1011011",
							neighbor35	WHEN "1011100",
							neighbor34	WHEN OTHERS;
							
	WITH mux_left SELECT
	neighbor_left1 <=	neighbor127	WHEN "0000000",
							neighbor126	WHEN "0000001",
							neighbor125	WHEN "0000010",
							neighbor124	WHEN "0000011",
							neighbor123	WHEN "0000100",
							neighbor122	WHEN "0000101",
							neighbor121	WHEN "0000110",
							neighbor120	WHEN "0000111",
							neighbor119	WHEN "0001000",
							neighbor118	WHEN "0001001",
							neighbor117	WHEN "0001010",
							neighbor116	WHEN "0001011",
							neighbor115	WHEN "0001100",
							neighbor114	WHEN "0001101",
							neighbor113	WHEN "0001110",
							neighbor112	WHEN "0001111",
							neighbor111	WHEN "0010000",
							neighbor110	WHEN "0010001",
							neighbor109	WHEN "0010010",
							neighbor108	WHEN "0010011",
							neighbor107	WHEN "0010100",
							neighbor106	WHEN "0010101",
							neighbor105	WHEN "0010110",
							neighbor104	WHEN "0010111",
							neighbor103	WHEN "0011000",
							neighbor102	WHEN "0011001",
							neighbor101	WHEN "0011010",
							neighbor100	WHEN "0011011",
							neighbor99	WHEN "0011100",
							neighbor98	WHEN "0011101",
							neighbor97	WHEN "0011110",
							neighbor96	WHEN "0011111",
							neighbor95	WHEN "0100000",
							neighbor94	WHEN "0100001",
							neighbor93	WHEN "0100010",
							neighbor92	WHEN "0100011",
							neighbor91	WHEN "0100100",
							neighbor90	WHEN "0100101",
							neighbor89	WHEN "0100110",
							neighbor88	WHEN "0100111",
							neighbor87	WHEN "0101000",
							neighbor86	WHEN "0101001",
							neighbor85	WHEN "0101010",
							neighbor84	WHEN "0101011",
							neighbor83	WHEN "0101100",
							neighbor82	WHEN "0101101",
							neighbor81	WHEN "0101110",
							neighbor80	WHEN "0101111",
							neighbor79	WHEN "0110000",
							neighbor78	WHEN "0110001",
							neighbor77	WHEN "0110010",
							neighbor76	WHEN "0110011",
							neighbor75	WHEN "0110100",
							neighbor74	WHEN "0110101",
							neighbor73	WHEN "0110110",
							neighbor72	WHEN "0110111",
							neighbor71	WHEN "0111000",
							neighbor70	WHEN "0111001",
							neighbor69	WHEN "0111010",
							neighbor68	WHEN "0111011",
							neighbor67	WHEN "0111100",
							neighbor66	WHEN "0111101",
							neighbor65	WHEN "0111110",
							neighborDC	WHEN "0111111",
							neighbor64	WHEN "1000000",
							neighbor63	WHEN "1000001",
							neighbor62	WHEN "1000010",
							neighbor61	WHEN "1000011",
							neighbor60	WHEN "1000100",
							neighbor59	WHEN "1000101",
							neighbor58	WHEN "1000110",
							neighbor57	WHEN "1000111",
							neighbor56	WHEN "1001000",
							neighbor55	WHEN "1001001",
							neighbor54	WHEN "1001010",
							neighbor53	WHEN "1001011",
							neighbor52	WHEN "1001100",
							neighbor51	WHEN "1001101",
							neighbor50	WHEN "1001110",
							neighbor49	WHEN "1001111",
							neighbor48	WHEN "1010000",
							neighbor47	WHEN "1010001",
							neighbor46	WHEN "1010010",
							neighbor45	WHEN "1010011",
							neighbor44	WHEN "1010100",
							neighbor43	WHEN "1010101",
							neighbor42	WHEN "1010110",
							neighbor41	WHEN "1010111",
							neighbor40	WHEN "1011000",
							neighbor39	WHEN "1011001",
							neighbor38	WHEN "1011010",
							neighbor37	WHEN "1011011",
							neighbor36	WHEN "1011100",
							neighbor35	WHEN OTHERS;
	
	WITH mux_left SELECT
	neighbor_left0 <=	neighbor127	WHEN "0000000",
							neighbor127	WHEN "0000001",
							neighbor126	WHEN "0000010",
							neighbor125	WHEN "0000011",
							neighbor124	WHEN "0000100",
							neighbor123	WHEN "0000101",
							neighbor122	WHEN "0000110",
							neighbor121	WHEN "0000111",
							neighbor120	WHEN "0001000",
							neighbor119	WHEN "0001001",
							neighbor118	WHEN "0001010",
							neighbor117	WHEN "0001011",
							neighbor116	WHEN "0001100",
							neighbor115	WHEN "0001101",
							neighbor114	WHEN "0001110",
							neighbor113	WHEN "0001111",
							neighbor112	WHEN "0010000",
							neighbor111	WHEN "0010001",
							neighbor110	WHEN "0010010",
							neighbor109	WHEN "0010011",
							neighbor108	WHEN "0010100",
							neighbor107	WHEN "0010101",
							neighbor106	WHEN "0010110",
							neighbor105	WHEN "0010111",
							neighbor104	WHEN "0011000",
							neighbor103	WHEN "0011001",
							neighbor102	WHEN "0011010",
							neighbor101	WHEN "0011011",
							neighbor100	WHEN "0011100",
							neighbor99	WHEN "0011101",
							neighbor98	WHEN "0011110",
							neighbor97	WHEN "0011111",
							neighbor96	WHEN "0100000",
							neighbor95	WHEN "0100001",
							neighbor94	WHEN "0100010",
							neighbor93	WHEN "0100011",
							neighbor92	WHEN "0100100",
							neighbor91	WHEN "0100101",
							neighbor90	WHEN "0100110",
							neighbor89	WHEN "0100111",
							neighbor88	WHEN "0101000",
							neighbor87	WHEN "0101001",
							neighbor86	WHEN "0101010",
							neighbor85	WHEN "0101011",
							neighbor84	WHEN "0101100",
							neighbor83	WHEN "0101101",
							neighbor82	WHEN "0101110",
							neighbor81	WHEN "0101111",
							neighbor80	WHEN "0110000",
							neighbor79	WHEN "0110001",
							neighbor78	WHEN "0110010",
							neighbor77	WHEN "0110011",
							neighbor76	WHEN "0110100",
							neighbor75	WHEN "0110101",
							neighbor74	WHEN "0110110",
							neighbor73	WHEN "0110111",
							neighbor72	WHEN "0111000",
							neighbor71	WHEN "0111001",
							neighbor70	WHEN "0111010",
							neighbor69	WHEN "0111011",
							neighbor68	WHEN "0111100",
							neighbor67	WHEN "0111101",
							neighbor66	WHEN "0111110",
							neighbor65	WHEN "0111111",
							neighborDC	WHEN "1000000",
							neighbor64	WHEN "1000001",
							neighbor63	WHEN "1000010",
							neighbor62	WHEN "1000011",
							neighbor61	WHEN "1000100",
							neighbor60	WHEN "1000101",
							neighbor59	WHEN "1000110",
							neighbor58	WHEN "1000111",
							neighbor57	WHEN "1001000",
							neighbor56	WHEN "1001001",
							neighbor55	WHEN "1001010",
							neighbor54	WHEN "1001011",
							neighbor53	WHEN "1001100",
							neighbor52	WHEN "1001101",
							neighbor51	WHEN "1001110",
							neighbor50	WHEN "1001111",
							neighbor49	WHEN "1010000",
							neighbor48	WHEN "1010001",
							neighbor47	WHEN "1010010",
							neighbor46	WHEN "1010011",
							neighbor45	WHEN "1010100",
							neighbor44	WHEN "1010101",
							neighbor43	WHEN "1010110",
							neighbor42	WHEN "1010111",
							neighbor41	WHEN "1011000",
							neighbor40	WHEN "1011001",
							neighbor39	WHEN "1011010",
							neighbor38	WHEN "1011011",
							neighbor37	WHEN "1011100",
							neighbor36	WHEN OTHERS;
							
END behavior;